---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
---------------------------------------------------------------------------
entity rom_img is

  port(addr : in  std_logic_vector(16 downto 0);
       clk  : in  std_logic;
       q    : out std_logic_vector(15 downto 0));

end entity;
---------------------------------------------------------------------------
architecture rtl of rom_img is

  -- Build a 2-D array type for the ROM
  subtype word_t is std_logic_vector(q'range);                 -- word size = q size
  type memory_t is array(0 to (2**addr'length) - 1) of word_t; -- number of words = 2^nbits(addr)

  function init_rom
    return memory_t is
    variable tmp : memory_t := (others => (others => '0'));
  begin
    tmp(00000) := x"0000";
    tmp(00001) := x"0020";
    tmp(00002) := x"0020";
    tmp(00003) := x"0020";
    tmp(00004) := x"0020";
    tmp(00005) := x"0020";
    tmp(00006) := x"0020";
    tmp(00007) := x"0020";
    tmp(00008) := x"0020";
    tmp(00009) := x"0020";
    tmp(00010) := x"0020";
    tmp(00011) := x"0020";
    tmp(00012) := x"0020";
    tmp(00013) := x"0020";
    tmp(00014) := x"0020";
    tmp(00015) := x"0040";
    tmp(00016) := x"0040";
    tmp(00017) := x"0040";
    tmp(00018) := x"0040";
    tmp(00019) := x"0040";
    tmp(00020) := x"0040";
    tmp(00021) := x"0060";
    tmp(00022) := x"0060";
    tmp(00023) := x"0860";
    tmp(00024) := x"0860";
    tmp(00025) := x"0860";
    tmp(00026) := x"0860";
    tmp(00027) := x"0860";
    tmp(00028) := x"0860";
    tmp(00029) := x"0860";
    tmp(00030) := x"0860";
    tmp(00031) := x"0060";
    tmp(00032) := x"0040";
    tmp(00033) := x"0040";
    tmp(00034) := x"0040";
    tmp(00035) := x"0040";
    tmp(00036) := x"0040";
    tmp(00037) := x"0040";
    tmp(00038) := x"0040";
    tmp(00039) := x"0040";
    tmp(00040) := x"0040";
    tmp(00041) := x"0040";
    tmp(00042) := x"0040";
    tmp(00043) := x"0040";
    tmp(00044) := x"0040";
    tmp(00045) := x"0020";
    tmp(00046) := x"0020";
    tmp(00047) := x"0020";
    tmp(00048) := x"0020";
    tmp(00049) := x"0020";
    tmp(00050) := x"0020";
    tmp(00051) := x"0020";
    tmp(00052) := x"0020";
    tmp(00053) := x"0020";
    tmp(00054) := x"0020";
    tmp(00055) := x"0020";
    tmp(00056) := x"0020";
    tmp(00057) := x"0020";
    tmp(00058) := x"0020";
    tmp(00059) := x"0040";
    tmp(00060) := x"0040";
    tmp(00061) := x"0040";
    tmp(00062) := x"0040";
    tmp(00063) := x"0040";
    tmp(00064) := x"0060";
    tmp(00065) := x"0060";
    tmp(00066) := x"0060";
    tmp(00067) := x"0860";
    tmp(00068) := x"0880";
    tmp(00069) := x"0880";
    tmp(00070) := x"0880";
    tmp(00071) := x"0880";
    tmp(00072) := x"08a0";
    tmp(00073) := x"08a0";
    tmp(00074) := x"08a0";
    tmp(00075) := x"08a0";
    tmp(00076) := x"08a0";
    tmp(00077) := x"08a0";
    tmp(00078) := x"08a0";
    tmp(00079) := x"08a0";
    tmp(00080) := x"08a0";
    tmp(00081) := x"08a0";
    tmp(00082) := x"08a0";
    tmp(00083) := x"08a0";
    tmp(00084) := x"08a0";
    tmp(00085) := x"08a0";
    tmp(00086) := x"08a0";
    tmp(00087) := x"08a0";
    tmp(00088) := x"08a0";
    tmp(00089) := x"08a0";
    tmp(00090) := x"08a0";
    tmp(00091) := x"08a0";
    tmp(00092) := x"08a0";
    tmp(00093) := x"08a0";
    tmp(00094) := x"08a0";
    tmp(00095) := x"08a0";
    tmp(00096) := x"08a0";
    tmp(00097) := x"08a0";
    tmp(00098) := x"08a0";
    tmp(00099) := x"08a0";
    tmp(00100) := x"08a0";
    tmp(00101) := x"08a0";
    tmp(00102) := x"08a0";
    tmp(00103) := x"08a0";
    tmp(00104) := x"08a0";
    tmp(00105) := x"08a0";
    tmp(00106) := x"08a0";
    tmp(00107) := x"08a0";
    tmp(00108) := x"08a0";
    tmp(00109) := x"08a0";
    tmp(00110) := x"08a0";
    tmp(00111) := x"08a0";
    tmp(00112) := x"08a0";
    tmp(00113) := x"08a0";
    tmp(00114) := x"08c0";
    tmp(00115) := x"08a0";
    tmp(00116) := x"08a0";
    tmp(00117) := x"08a0";
    tmp(00118) := x"08c0";
    tmp(00119) := x"08c0";
    tmp(00120) := x"08a0";
    tmp(00121) := x"08a0";
    tmp(00122) := x"08a0";
    tmp(00123) := x"08a0";
    tmp(00124) := x"08a0";
    tmp(00125) := x"08a0";
    tmp(00126) := x"08a0";
    tmp(00127) := x"08a0";
    tmp(00128) := x"08a0";
    tmp(00129) := x"08a0";
    tmp(00130) := x"08a0";
    tmp(00131) := x"08a0";
    tmp(00132) := x"08a0";
    tmp(00133) := x"08a0";
    tmp(00134) := x"08a0";
    tmp(00135) := x"08a0";
    tmp(00136) := x"08a0";
    tmp(00137) := x"08a0";
    tmp(00138) := x"08a0";
    tmp(00139) := x"08a0";
    tmp(00140) := x"08a0";
    tmp(00141) := x"08a0";
    tmp(00142) := x"08a0";
    tmp(00143) := x"08a0";
    tmp(00144) := x"08a0";
    tmp(00145) := x"08a0";
    tmp(00146) := x"08a0";
    tmp(00147) := x"08a0";
    tmp(00148) := x"08a0";
    tmp(00149) := x"08a0";
    tmp(00150) := x"08a0";
    tmp(00151) := x"08a0";
    tmp(00152) := x"08a0";
    tmp(00153) := x"08a0";
    tmp(00154) := x"08a0";
    tmp(00155) := x"08a0";
    tmp(00156) := x"08a0";
    tmp(00157) := x"08a0";
    tmp(00158) := x"08a0";
    tmp(00159) := x"08a0";
    tmp(00160) := x"08a0";
    tmp(00161) := x"08a0";
    tmp(00162) := x"08a0";
    tmp(00163) := x"08a0";
    tmp(00164) := x"08a0";
    tmp(00165) := x"08a0";
    tmp(00166) := x"08a0";
    tmp(00167) := x"08a0";
    tmp(00168) := x"08a0";
    tmp(00169) := x"08a0";
    tmp(00170) := x"08a0";
    tmp(00171) := x"08a0";
    tmp(00172) := x"08a0";
    tmp(00173) := x"08a0";
    tmp(00174) := x"08a0";
    tmp(00175) := x"08a0";
    tmp(00176) := x"08a0";
    tmp(00177) := x"08a0";
    tmp(00178) := x"08a0";
    tmp(00179) := x"08a0";
    tmp(00180) := x"08a0";
    tmp(00181) := x"08a0";
    tmp(00182) := x"08a0";
    tmp(00183) := x"08a0";
    tmp(00184) := x"08a0";
    tmp(00185) := x"08a0";
    tmp(00186) := x"08a0";
    tmp(00187) := x"08a0";
    tmp(00188) := x"08a0";
    tmp(00189) := x"08a0";
    tmp(00190) := x"08a0";
    tmp(00191) := x"08a0";
    tmp(00192) := x"08a0";
    tmp(00193) := x"08a0";
    tmp(00194) := x"08a0";
    tmp(00195) := x"08a0";
    tmp(00196) := x"08a0";
    tmp(00197) := x"08a0";
    tmp(00198) := x"08a0";
    tmp(00199) := x"08a0";
    tmp(00200) := x"08a0";
    tmp(00201) := x"08a0";
    tmp(00202) := x"08a0";
    tmp(00203) := x"0880";
    tmp(00204) := x"0880";
    tmp(00205) := x"0880";
    tmp(00206) := x"0880";
    tmp(00207) := x"0880";
    tmp(00208) := x"0880";
    tmp(00209) := x"0880";
    tmp(00210) := x"0880";
    tmp(00211) := x"0880";
    tmp(00212) := x"0880";
    tmp(00213) := x"0880";
    tmp(00214) := x"0860";
    tmp(00215) := x"0860";
    tmp(00216) := x"0860";
    tmp(00217) := x"0860";
    tmp(00218) := x"0860";
    tmp(00219) := x"0860";
    tmp(00220) := x"0860";
    tmp(00221) := x"0860";
    tmp(00222) := x"0840";
    tmp(00223) := x"0840";
    tmp(00224) := x"0840";
    tmp(00225) := x"0840";
    tmp(00226) := x"0840";
    tmp(00227) := x"0840";
    tmp(00228) := x"0840";
    tmp(00229) := x"0820";
    tmp(00230) := x"0820";
    tmp(00231) := x"0820";
    tmp(00232) := x"0820";
    tmp(00233) := x"0820";
    tmp(00234) := x"0820";
    tmp(00235) := x"0820";
    tmp(00236) := x"0820";
    tmp(00237) := x"0820";
    tmp(00238) := x"0820";
    tmp(00239) := x"0820";
    tmp(00240) := x"0000";
    tmp(00241) := x"0020";
    tmp(00242) := x"0020";
    tmp(00243) := x"0020";
    tmp(00244) := x"0020";
    tmp(00245) := x"0020";
    tmp(00246) := x"0020";
    tmp(00247) := x"0020";
    tmp(00248) := x"0020";
    tmp(00249) := x"0020";
    tmp(00250) := x"0020";
    tmp(00251) := x"0020";
    tmp(00252) := x"0020";
    tmp(00253) := x"0020";
    tmp(00254) := x"0020";
    tmp(00255) := x"0020";
    tmp(00256) := x"0040";
    tmp(00257) := x"0040";
    tmp(00258) := x"0040";
    tmp(00259) := x"0040";
    tmp(00260) := x"0040";
    tmp(00261) := x"0040";
    tmp(00262) := x"0060";
    tmp(00263) := x"0860";
    tmp(00264) := x"0860";
    tmp(00265) := x"0860";
    tmp(00266) := x"0860";
    tmp(00267) := x"0860";
    tmp(00268) := x"0860";
    tmp(00269) := x"0860";
    tmp(00270) := x"0860";
    tmp(00271) := x"0860";
    tmp(00272) := x"0040";
    tmp(00273) := x"0040";
    tmp(00274) := x"0040";
    tmp(00275) := x"0040";
    tmp(00276) := x"0040";
    tmp(00277) := x"0040";
    tmp(00278) := x"0040";
    tmp(00279) := x"0040";
    tmp(00280) := x"0040";
    tmp(00281) := x"0040";
    tmp(00282) := x"0040";
    tmp(00283) := x"0040";
    tmp(00284) := x"0020";
    tmp(00285) := x"0020";
    tmp(00286) := x"0020";
    tmp(00287) := x"0020";
    tmp(00288) := x"0020";
    tmp(00289) := x"0020";
    tmp(00290) := x"0020";
    tmp(00291) := x"0020";
    tmp(00292) := x"0020";
    tmp(00293) := x"0020";
    tmp(00294) := x"0020";
    tmp(00295) := x"0020";
    tmp(00296) := x"0040";
    tmp(00297) := x"0040";
    tmp(00298) := x"0040";
    tmp(00299) := x"0040";
    tmp(00300) := x"0040";
    tmp(00301) := x"0040";
    tmp(00302) := x"0060";
    tmp(00303) := x"0060";
    tmp(00304) := x"0060";
    tmp(00305) := x"0880";
    tmp(00306) := x"0880";
    tmp(00307) := x"0880";
    tmp(00308) := x"0880";
    tmp(00309) := x"0880";
    tmp(00310) := x"08a0";
    tmp(00311) := x"08a0";
    tmp(00312) := x"08a0";
    tmp(00313) := x"08a0";
    tmp(00314) := x"08a0";
    tmp(00315) := x"08a0";
    tmp(00316) := x"08a0";
    tmp(00317) := x"08a0";
    tmp(00318) := x"08a0";
    tmp(00319) := x"08a0";
    tmp(00320) := x"08a0";
    tmp(00321) := x"0880";
    tmp(00322) := x"08a0";
    tmp(00323) := x"0880";
    tmp(00324) := x"0880";
    tmp(00325) := x"0880";
    tmp(00326) := x"0880";
    tmp(00327) := x"0880";
    tmp(00328) := x"0880";
    tmp(00329) := x"08a0";
    tmp(00330) := x"0880";
    tmp(00331) := x"08a0";
    tmp(00332) := x"08a0";
    tmp(00333) := x"08a0";
    tmp(00334) := x"08a0";
    tmp(00335) := x"0880";
    tmp(00336) := x"08a0";
    tmp(00337) := x"08a0";
    tmp(00338) := x"08a0";
    tmp(00339) := x"08a0";
    tmp(00340) := x"0880";
    tmp(00341) := x"0880";
    tmp(00342) := x"0880";
    tmp(00343) := x"0880";
    tmp(00344) := x"0880";
    tmp(00345) := x"0880";
    tmp(00346) := x"08a0";
    tmp(00347) := x"08a0";
    tmp(00348) := x"0880";
    tmp(00349) := x"08a0";
    tmp(00350) := x"08a0";
    tmp(00351) := x"08a0";
    tmp(00352) := x"08a0";
    tmp(00353) := x"08a0";
    tmp(00354) := x"08a0";
    tmp(00355) := x"08a0";
    tmp(00356) := x"08a0";
    tmp(00357) := x"08a0";
    tmp(00358) := x"08a0";
    tmp(00359) := x"08a0";
    tmp(00360) := x"08a0";
    tmp(00361) := x"08a0";
    tmp(00362) := x"08a0";
    tmp(00363) := x"08a0";
    tmp(00364) := x"08a0";
    tmp(00365) := x"08a0";
    tmp(00366) := x"08a0";
    tmp(00367) := x"08a0";
    tmp(00368) := x"08a0";
    tmp(00369) := x"08a0";
    tmp(00370) := x"08a0";
    tmp(00371) := x"08a0";
    tmp(00372) := x"08a0";
    tmp(00373) := x"08a0";
    tmp(00374) := x"08a0";
    tmp(00375) := x"08a0";
    tmp(00376) := x"08a0";
    tmp(00377) := x"08a0";
    tmp(00378) := x"08a0";
    tmp(00379) := x"08a0";
    tmp(00380) := x"08a0";
    tmp(00381) := x"08a0";
    tmp(00382) := x"08a0";
    tmp(00383) := x"08a0";
    tmp(00384) := x"08a0";
    tmp(00385) := x"08a0";
    tmp(00386) := x"08a0";
    tmp(00387) := x"08a0";
    tmp(00388) := x"08a0";
    tmp(00389) := x"08a0";
    tmp(00390) := x"08a0";
    tmp(00391) := x"08a0";
    tmp(00392) := x"08a0";
    tmp(00393) := x"08a0";
    tmp(00394) := x"08a0";
    tmp(00395) := x"08a0";
    tmp(00396) := x"08a0";
    tmp(00397) := x"08a0";
    tmp(00398) := x"08a0";
    tmp(00399) := x"08a0";
    tmp(00400) := x"0880";
    tmp(00401) := x"08a0";
    tmp(00402) := x"08a0";
    tmp(00403) := x"08a0";
    tmp(00404) := x"08a0";
    tmp(00405) := x"08a0";
    tmp(00406) := x"08a0";
    tmp(00407) := x"0880";
    tmp(00408) := x"0880";
    tmp(00409) := x"08a0";
    tmp(00410) := x"0880";
    tmp(00411) := x"0880";
    tmp(00412) := x"0880";
    tmp(00413) := x"08a0";
    tmp(00414) := x"08a0";
    tmp(00415) := x"08a0";
    tmp(00416) := x"08a0";
    tmp(00417) := x"08a0";
    tmp(00418) := x"08a0";
    tmp(00419) := x"08a0";
    tmp(00420) := x"08a0";
    tmp(00421) := x"08a0";
    tmp(00422) := x"08a0";
    tmp(00423) := x"08a0";
    tmp(00424) := x"08a0";
    tmp(00425) := x"08a0";
    tmp(00426) := x"08a0";
    tmp(00427) := x"08a0";
    tmp(00428) := x"08a0";
    tmp(00429) := x"08a0";
    tmp(00430) := x"08a0";
    tmp(00431) := x"08a0";
    tmp(00432) := x"08a0";
    tmp(00433) := x"08a0";
    tmp(00434) := x"08a0";
    tmp(00435) := x"08a0";
    tmp(00436) := x"08a0";
    tmp(00437) := x"08a0";
    tmp(00438) := x"08a0";
    tmp(00439) := x"08a0";
    tmp(00440) := x"08a0";
    tmp(00441) := x"08a0";
    tmp(00442) := x"0880";
    tmp(00443) := x"0880";
    tmp(00444) := x"0880";
    tmp(00445) := x"0880";
    tmp(00446) := x"0880";
    tmp(00447) := x"0880";
    tmp(00448) := x"0880";
    tmp(00449) := x"0880";
    tmp(00450) := x"0880";
    tmp(00451) := x"0860";
    tmp(00452) := x"0860";
    tmp(00453) := x"0860";
    tmp(00454) := x"0860";
    tmp(00455) := x"0860";
    tmp(00456) := x"0860";
    tmp(00457) := x"0860";
    tmp(00458) := x"0860";
    tmp(00459) := x"0860";
    tmp(00460) := x"0860";
    tmp(00461) := x"0860";
    tmp(00462) := x"0860";
    tmp(00463) := x"0840";
    tmp(00464) := x"0840";
    tmp(00465) := x"0840";
    tmp(00466) := x"0840";
    tmp(00467) := x"0840";
    tmp(00468) := x"0840";
    tmp(00469) := x"0820";
    tmp(00470) := x"0820";
    tmp(00471) := x"0820";
    tmp(00472) := x"0820";
    tmp(00473) := x"0820";
    tmp(00474) := x"0820";
    tmp(00475) := x"0820";
    tmp(00476) := x"0820";
    tmp(00477) := x"0820";
    tmp(00478) := x"0820";
    tmp(00479) := x"0820";
    tmp(00480) := x"0000";
    tmp(00481) := x"0020";
    tmp(00482) := x"0000";
    tmp(00483) := x"0020";
    tmp(00484) := x"0020";
    tmp(00485) := x"0020";
    tmp(00486) := x"0020";
    tmp(00487) := x"0020";
    tmp(00488) := x"0020";
    tmp(00489) := x"0020";
    tmp(00490) := x"0020";
    tmp(00491) := x"0020";
    tmp(00492) := x"0020";
    tmp(00493) := x"0020";
    tmp(00494) := x"0020";
    tmp(00495) := x"0020";
    tmp(00496) := x"0020";
    tmp(00497) := x"0040";
    tmp(00498) := x"0040";
    tmp(00499) := x"0040";
    tmp(00500) := x"0040";
    tmp(00501) := x"0040";
    tmp(00502) := x"0060";
    tmp(00503) := x"0860";
    tmp(00504) := x"0860";
    tmp(00505) := x"0860";
    tmp(00506) := x"0860";
    tmp(00507) := x"0860";
    tmp(00508) := x"0860";
    tmp(00509) := x"0860";
    tmp(00510) := x"0060";
    tmp(00511) := x"0040";
    tmp(00512) := x"0040";
    tmp(00513) := x"0040";
    tmp(00514) := x"0040";
    tmp(00515) := x"0040";
    tmp(00516) := x"0040";
    tmp(00517) := x"0040";
    tmp(00518) := x"0040";
    tmp(00519) := x"0040";
    tmp(00520) := x"0040";
    tmp(00521) := x"0040";
    tmp(00522) := x"0040";
    tmp(00523) := x"0020";
    tmp(00524) := x"0020";
    tmp(00525) := x"0020";
    tmp(00526) := x"0020";
    tmp(00527) := x"0020";
    tmp(00528) := x"0020";
    tmp(00529) := x"0020";
    tmp(00530) := x"0020";
    tmp(00531) := x"0020";
    tmp(00532) := x"0020";
    tmp(00533) := x"0020";
    tmp(00534) := x"0040";
    tmp(00535) := x"0040";
    tmp(00536) := x"0040";
    tmp(00537) := x"0040";
    tmp(00538) := x"0040";
    tmp(00539) := x"0040";
    tmp(00540) := x"0060";
    tmp(00541) := x"0060";
    tmp(00542) := x"0860";
    tmp(00543) := x"0860";
    tmp(00544) := x"0880";
    tmp(00545) := x"0880";
    tmp(00546) := x"0880";
    tmp(00547) := x"0880";
    tmp(00548) := x"08a0";
    tmp(00549) := x"08a0";
    tmp(00550) := x"08a0";
    tmp(00551) := x"08a0";
    tmp(00552) := x"08a0";
    tmp(00553) := x"08a0";
    tmp(00554) := x"08a0";
    tmp(00555) := x"08a0";
    tmp(00556) := x"08a0";
    tmp(00557) := x"08a0";
    tmp(00558) := x"0880";
    tmp(00559) := x"0880";
    tmp(00560) := x"0880";
    tmp(00561) := x"0880";
    tmp(00562) := x"0880";
    tmp(00563) := x"0880";
    tmp(00564) := x"0880";
    tmp(00565) := x"0880";
    tmp(00566) := x"0880";
    tmp(00567) := x"0880";
    tmp(00568) := x"0880";
    tmp(00569) := x"0880";
    tmp(00570) := x"0880";
    tmp(00571) := x"0880";
    tmp(00572) := x"0880";
    tmp(00573) := x"0880";
    tmp(00574) := x"0880";
    tmp(00575) := x"0880";
    tmp(00576) := x"0880";
    tmp(00577) := x"0880";
    tmp(00578) := x"0880";
    tmp(00579) := x"0880";
    tmp(00580) := x"0880";
    tmp(00581) := x"0880";
    tmp(00582) := x"0880";
    tmp(00583) := x"0880";
    tmp(00584) := x"0880";
    tmp(00585) := x"0880";
    tmp(00586) := x"0880";
    tmp(00587) := x"0880";
    tmp(00588) := x"0880";
    tmp(00589) := x"0880";
    tmp(00590) := x"08a0";
    tmp(00591) := x"08a0";
    tmp(00592) := x"08a0";
    tmp(00593) := x"08a0";
    tmp(00594) := x"08a0";
    tmp(00595) := x"08a0";
    tmp(00596) := x"08a0";
    tmp(00597) := x"08a0";
    tmp(00598) := x"08a0";
    tmp(00599) := x"08a0";
    tmp(00600) := x"08a0";
    tmp(00601) := x"08a0";
    tmp(00602) := x"08a0";
    tmp(00603) := x"08a0";
    tmp(00604) := x"08a0";
    tmp(00605) := x"08a0";
    tmp(00606) := x"08a0";
    tmp(00607) := x"08a0";
    tmp(00608) := x"08a0";
    tmp(00609) := x"08a0";
    tmp(00610) := x"08a0";
    tmp(00611) := x"08a0";
    tmp(00612) := x"08a0";
    tmp(00613) := x"08a0";
    tmp(00614) := x"08a0";
    tmp(00615) := x"08a0";
    tmp(00616) := x"08a0";
    tmp(00617) := x"08a0";
    tmp(00618) := x"08a0";
    tmp(00619) := x"08a0";
    tmp(00620) := x"08a0";
    tmp(00621) := x"08a0";
    tmp(00622) := x"08a0";
    tmp(00623) := x"08a0";
    tmp(00624) := x"08a0";
    tmp(00625) := x"08a0";
    tmp(00626) := x"08a0";
    tmp(00627) := x"08a0";
    tmp(00628) := x"08a0";
    tmp(00629) := x"08a0";
    tmp(00630) := x"08a0";
    tmp(00631) := x"08a0";
    tmp(00632) := x"08a0";
    tmp(00633) := x"08a0";
    tmp(00634) := x"08a0";
    tmp(00635) := x"08a0";
    tmp(00636) := x"08a0";
    tmp(00637) := x"08a0";
    tmp(00638) := x"08a0";
    tmp(00639) := x"08a0";
    tmp(00640) := x"08a0";
    tmp(00641) := x"08a0";
    tmp(00642) := x"08a0";
    tmp(00643) := x"08a0";
    tmp(00644) := x"08a0";
    tmp(00645) := x"08a0";
    tmp(00646) := x"0880";
    tmp(00647) := x"0880";
    tmp(00648) := x"0880";
    tmp(00649) := x"0880";
    tmp(00650) := x"0880";
    tmp(00651) := x"0880";
    tmp(00652) := x"0880";
    tmp(00653) := x"0880";
    tmp(00654) := x"0880";
    tmp(00655) := x"0880";
    tmp(00656) := x"0880";
    tmp(00657) := x"0880";
    tmp(00658) := x"0880";
    tmp(00659) := x"0880";
    tmp(00660) := x"0880";
    tmp(00661) := x"0880";
    tmp(00662) := x"08a0";
    tmp(00663) := x"08a0";
    tmp(00664) := x"0880";
    tmp(00665) := x"0880";
    tmp(00666) := x"08a0";
    tmp(00667) := x"08a0";
    tmp(00668) := x"08a0";
    tmp(00669) := x"08a0";
    tmp(00670) := x"08a0";
    tmp(00671) := x"08a0";
    tmp(00672) := x"08a0";
    tmp(00673) := x"08a0";
    tmp(00674) := x"08a0";
    tmp(00675) := x"08a0";
    tmp(00676) := x"08a0";
    tmp(00677) := x"08a0";
    tmp(00678) := x"08a0";
    tmp(00679) := x"08a0";
    tmp(00680) := x"08a0";
    tmp(00681) := x"0880";
    tmp(00682) := x"0880";
    tmp(00683) := x"0880";
    tmp(00684) := x"0880";
    tmp(00685) := x"0880";
    tmp(00686) := x"0880";
    tmp(00687) := x"0880";
    tmp(00688) := x"0880";
    tmp(00689) := x"0880";
    tmp(00690) := x"0860";
    tmp(00691) := x"0860";
    tmp(00692) := x"0860";
    tmp(00693) := x"0860";
    tmp(00694) := x"0860";
    tmp(00695) := x"0860";
    tmp(00696) := x"0860";
    tmp(00697) := x"0860";
    tmp(00698) := x"0860";
    tmp(00699) := x"0860";
    tmp(00700) := x"0860";
    tmp(00701) := x"0860";
    tmp(00702) := x"0860";
    tmp(00703) := x"0840";
    tmp(00704) := x"0840";
    tmp(00705) := x"0840";
    tmp(00706) := x"0840";
    tmp(00707) := x"0840";
    tmp(00708) := x"0840";
    tmp(00709) := x"0820";
    tmp(00710) := x"0820";
    tmp(00711) := x"0820";
    tmp(00712) := x"0820";
    tmp(00713) := x"0820";
    tmp(00714) := x"0820";
    tmp(00715) := x"0820";
    tmp(00716) := x"0820";
    tmp(00717) := x"0820";
    tmp(00718) := x"0820";
    tmp(00719) := x"0820";
    tmp(00720) := x"0000";
    tmp(00721) := x"0020";
    tmp(00722) := x"0020";
    tmp(00723) := x"0020";
    tmp(00724) := x"0020";
    tmp(00725) := x"0020";
    tmp(00726) := x"0020";
    tmp(00727) := x"0020";
    tmp(00728) := x"0020";
    tmp(00729) := x"0020";
    tmp(00730) := x"0020";
    tmp(00731) := x"0020";
    tmp(00732) := x"0020";
    tmp(00733) := x"0020";
    tmp(00734) := x"0020";
    tmp(00735) := x"0020";
    tmp(00736) := x"0040";
    tmp(00737) := x"0040";
    tmp(00738) := x"0040";
    tmp(00739) := x"0040";
    tmp(00740) := x"0040";
    tmp(00741) := x"0040";
    tmp(00742) := x"0060";
    tmp(00743) := x"0060";
    tmp(00744) := x"0060";
    tmp(00745) := x"0040";
    tmp(00746) := x"0040";
    tmp(00747) := x"0040";
    tmp(00748) := x"0040";
    tmp(00749) := x"0040";
    tmp(00750) := x"0040";
    tmp(00751) := x"0040";
    tmp(00752) := x"0040";
    tmp(00753) := x"0040";
    tmp(00754) := x"0040";
    tmp(00755) := x"0040";
    tmp(00756) := x"0040";
    tmp(00757) := x"0040";
    tmp(00758) := x"0040";
    tmp(00759) := x"0040";
    tmp(00760) := x"0040";
    tmp(00761) := x"0040";
    tmp(00762) := x"0020";
    tmp(00763) := x"0020";
    tmp(00764) := x"0020";
    tmp(00765) := x"0020";
    tmp(00766) := x"0020";
    tmp(00767) := x"0020";
    tmp(00768) := x"0020";
    tmp(00769) := x"0020";
    tmp(00770) := x"0020";
    tmp(00771) := x"0020";
    tmp(00772) := x"0040";
    tmp(00773) := x"0040";
    tmp(00774) := x"0040";
    tmp(00775) := x"0040";
    tmp(00776) := x"0040";
    tmp(00777) := x"0040";
    tmp(00778) := x"0060";
    tmp(00779) := x"0060";
    tmp(00780) := x"0060";
    tmp(00781) := x"0060";
    tmp(00782) := x"0860";
    tmp(00783) := x"0880";
    tmp(00784) := x"0880";
    tmp(00785) := x"0880";
    tmp(00786) := x"08a0";
    tmp(00787) := x"08a0";
    tmp(00788) := x"08a0";
    tmp(00789) := x"08a0";
    tmp(00790) := x"08a0";
    tmp(00791) := x"08a0";
    tmp(00792) := x"08a0";
    tmp(00793) := x"08a0";
    tmp(00794) := x"08a0";
    tmp(00795) := x"08a0";
    tmp(00796) := x"08a0";
    tmp(00797) := x"0880";
    tmp(00798) := x"0880";
    tmp(00799) := x"0880";
    tmp(00800) := x"0880";
    tmp(00801) := x"0880";
    tmp(00802) := x"0880";
    tmp(00803) := x"0880";
    tmp(00804) := x"0880";
    tmp(00805) := x"0880";
    tmp(00806) := x"0880";
    tmp(00807) := x"0880";
    tmp(00808) := x"0880";
    tmp(00809) := x"0880";
    tmp(00810) := x"0880";
    tmp(00811) := x"0880";
    tmp(00812) := x"0880";
    tmp(00813) := x"0880";
    tmp(00814) := x"0880";
    tmp(00815) := x"0880";
    tmp(00816) := x"0880";
    tmp(00817) := x"0880";
    tmp(00818) := x"0880";
    tmp(00819) := x"0880";
    tmp(00820) := x"0880";
    tmp(00821) := x"0880";
    tmp(00822) := x"0860";
    tmp(00823) := x"0860";
    tmp(00824) := x"0060";
    tmp(00825) := x"0060";
    tmp(00826) := x"0060";
    tmp(00827) := x"0060";
    tmp(00828) := x"0080";
    tmp(00829) := x"0080";
    tmp(00830) := x"0080";
    tmp(00831) := x"0880";
    tmp(00832) := x"0880";
    tmp(00833) := x"0880";
    tmp(00834) := x"0880";
    tmp(00835) := x"0880";
    tmp(00836) := x"08a0";
    tmp(00837) := x"0880";
    tmp(00838) := x"08a0";
    tmp(00839) := x"08a0";
    tmp(00840) := x"08a0";
    tmp(00841) := x"08a0";
    tmp(00842) := x"08a0";
    tmp(00843) := x"08a0";
    tmp(00844) := x"08a0";
    tmp(00845) := x"08a0";
    tmp(00846) := x"08a0";
    tmp(00847) := x"08a0";
    tmp(00848) := x"08a0";
    tmp(00849) := x"08a0";
    tmp(00850) := x"08a0";
    tmp(00851) := x"08a0";
    tmp(00852) := x"08a0";
    tmp(00853) := x"08a0";
    tmp(00854) := x"08a0";
    tmp(00855) := x"08a0";
    tmp(00856) := x"08a0";
    tmp(00857) := x"08a0";
    tmp(00858) := x"08a0";
    tmp(00859) := x"08a0";
    tmp(00860) := x"08a0";
    tmp(00861) := x"08a0";
    tmp(00862) := x"08a0";
    tmp(00863) := x"08a0";
    tmp(00864) := x"08a0";
    tmp(00865) := x"08a0";
    tmp(00866) := x"08a0";
    tmp(00867) := x"08a0";
    tmp(00868) := x"08a0";
    tmp(00869) := x"08a0";
    tmp(00870) := x"08a0";
    tmp(00871) := x"08a0";
    tmp(00872) := x"08a0";
    tmp(00873) := x"08a0";
    tmp(00874) := x"08a0";
    tmp(00875) := x"08a0";
    tmp(00876) := x"08a0";
    tmp(00877) := x"08a0";
    tmp(00878) := x"08a0";
    tmp(00879) := x"08a0";
    tmp(00880) := x"08a0";
    tmp(00881) := x"08a0";
    tmp(00882) := x"08a0";
    tmp(00883) := x"08a0";
    tmp(00884) := x"08a0";
    tmp(00885) := x"08a0";
    tmp(00886) := x"08a0";
    tmp(00887) := x"0880";
    tmp(00888) := x"0880";
    tmp(00889) := x"0880";
    tmp(00890) := x"0880";
    tmp(00891) := x"0880";
    tmp(00892) := x"0880";
    tmp(00893) := x"0880";
    tmp(00894) := x"0880";
    tmp(00895) := x"0880";
    tmp(00896) := x"0880";
    tmp(00897) := x"0880";
    tmp(00898) := x"0880";
    tmp(00899) := x"0880";
    tmp(00900) := x"0880";
    tmp(00901) := x"0880";
    tmp(00902) := x"0880";
    tmp(00903) := x"0880";
    tmp(00904) := x"0880";
    tmp(00905) := x"0880";
    tmp(00906) := x"0880";
    tmp(00907) := x"0880";
    tmp(00908) := x"0880";
    tmp(00909) := x"0880";
    tmp(00910) := x"0880";
    tmp(00911) := x"0880";
    tmp(00912) := x"0880";
    tmp(00913) := x"0880";
    tmp(00914) := x"0880";
    tmp(00915) := x"0880";
    tmp(00916) := x"0880";
    tmp(00917) := x"0880";
    tmp(00918) := x"0880";
    tmp(00919) := x"0880";
    tmp(00920) := x"0880";
    tmp(00921) := x"0880";
    tmp(00922) := x"0880";
    tmp(00923) := x"0880";
    tmp(00924) := x"0880";
    tmp(00925) := x"0880";
    tmp(00926) := x"0880";
    tmp(00927) := x"0880";
    tmp(00928) := x"0880";
    tmp(00929) := x"0880";
    tmp(00930) := x"0860";
    tmp(00931) := x"0860";
    tmp(00932) := x"0860";
    tmp(00933) := x"0860";
    tmp(00934) := x"0860";
    tmp(00935) := x"0860";
    tmp(00936) := x"0860";
    tmp(00937) := x"0860";
    tmp(00938) := x"0860";
    tmp(00939) := x"0860";
    tmp(00940) := x"0840";
    tmp(00941) := x"0840";
    tmp(00942) := x"0840";
    tmp(00943) := x"0840";
    tmp(00944) := x"0840";
    tmp(00945) := x"0840";
    tmp(00946) := x"0840";
    tmp(00947) := x"0840";
    tmp(00948) := x"0840";
    tmp(00949) := x"0840";
    tmp(00950) := x"0820";
    tmp(00951) := x"0820";
    tmp(00952) := x"0820";
    tmp(00953) := x"0820";
    tmp(00954) := x"0820";
    tmp(00955) := x"0820";
    tmp(00956) := x"0820";
    tmp(00957) := x"0820";
    tmp(00958) := x"0820";
    tmp(00959) := x"0820";
    tmp(00960) := x"0000";
    tmp(00961) := x"0020";
    tmp(00962) := x"0020";
    tmp(00963) := x"0020";
    tmp(00964) := x"0020";
    tmp(00965) := x"0020";
    tmp(00966) := x"0020";
    tmp(00967) := x"0020";
    tmp(00968) := x"0020";
    tmp(00969) := x"0020";
    tmp(00970) := x"0020";
    tmp(00971) := x"0020";
    tmp(00972) := x"0020";
    tmp(00973) := x"0020";
    tmp(00974) := x"0020";
    tmp(00975) := x"0020";
    tmp(00976) := x"0040";
    tmp(00977) := x"0040";
    tmp(00978) := x"0040";
    tmp(00979) := x"0040";
    tmp(00980) := x"0040";
    tmp(00981) := x"0040";
    tmp(00982) := x"0040";
    tmp(00983) := x"0040";
    tmp(00984) := x"0040";
    tmp(00985) := x"0040";
    tmp(00986) := x"0040";
    tmp(00987) := x"0040";
    tmp(00988) := x"0040";
    tmp(00989) := x"0040";
    tmp(00990) := x"0040";
    tmp(00991) := x"0040";
    tmp(00992) := x"0040";
    tmp(00993) := x"0040";
    tmp(00994) := x"0040";
    tmp(00995) := x"0040";
    tmp(00996) := x"0040";
    tmp(00997) := x"0040";
    tmp(00998) := x"0040";
    tmp(00999) := x"0040";
    tmp(01000) := x"0040";
    tmp(01001) := x"0040";
    tmp(01002) := x"0020";
    tmp(01003) := x"0020";
    tmp(01004) := x"0020";
    tmp(01005) := x"0040";
    tmp(01006) := x"0040";
    tmp(01007) := x"0040";
    tmp(01008) := x"0040";
    tmp(01009) := x"0040";
    tmp(01010) := x"0040";
    tmp(01011) := x"0040";
    tmp(01012) := x"0040";
    tmp(01013) := x"0040";
    tmp(01014) := x"0040";
    tmp(01015) := x"0040";
    tmp(01016) := x"0060";
    tmp(01017) := x"0060";
    tmp(01018) := x"0060";
    tmp(01019) := x"0060";
    tmp(01020) := x"0080";
    tmp(01021) := x"0880";
    tmp(01022) := x"0880";
    tmp(01023) := x"0880";
    tmp(01024) := x"0880";
    tmp(01025) := x"08a0";
    tmp(01026) := x"08a0";
    tmp(01027) := x"08a0";
    tmp(01028) := x"08a0";
    tmp(01029) := x"08a0";
    tmp(01030) := x"08a0";
    tmp(01031) := x"08a0";
    tmp(01032) := x"08a0";
    tmp(01033) := x"0880";
    tmp(01034) := x"0880";
    tmp(01035) := x"0880";
    tmp(01036) := x"0880";
    tmp(01037) := x"0880";
    tmp(01038) := x"0880";
    tmp(01039) := x"0880";
    tmp(01040) := x"0860";
    tmp(01041) := x"0860";
    tmp(01042) := x"0860";
    tmp(01043) := x"0860";
    tmp(01044) := x"0860";
    tmp(01045) := x"0860";
    tmp(01046) := x"0860";
    tmp(01047) := x"0860";
    tmp(01048) := x"0880";
    tmp(01049) := x"0880";
    tmp(01050) := x"0880";
    tmp(01051) := x"0880";
    tmp(01052) := x"0880";
    tmp(01053) := x"0880";
    tmp(01054) := x"0880";
    tmp(01055) := x"0880";
    tmp(01056) := x"0880";
    tmp(01057) := x"0880";
    tmp(01058) := x"0880";
    tmp(01059) := x"0880";
    tmp(01060) := x"0880";
    tmp(01061) := x"0860";
    tmp(01062) := x"0060";
    tmp(01063) := x"0060";
    tmp(01064) := x"0060";
    tmp(01065) := x"0060";
    tmp(01066) := x"0060";
    tmp(01067) := x"0060";
    tmp(01068) := x"0060";
    tmp(01069) := x"0060";
    tmp(01070) := x"0060";
    tmp(01071) := x"0060";
    tmp(01072) := x"0080";
    tmp(01073) := x"0080";
    tmp(01074) := x"0080";
    tmp(01075) := x"0080";
    tmp(01076) := x"0080";
    tmp(01077) := x"0080";
    tmp(01078) := x"0080";
    tmp(01079) := x"0080";
    tmp(01080) := x"0080";
    tmp(01081) := x"00a0";
    tmp(01082) := x"0080";
    tmp(01083) := x"00a0";
    tmp(01084) := x"00a0";
    tmp(01085) := x"00a0";
    tmp(01086) := x"00a0";
    tmp(01087) := x"08a0";
    tmp(01088) := x"08a0";
    tmp(01089) := x"08a0";
    tmp(01090) := x"08a0";
    tmp(01091) := x"08a0";
    tmp(01092) := x"08a0";
    tmp(01093) := x"08a0";
    tmp(01094) := x"08a0";
    tmp(01095) := x"08a0";
    tmp(01096) := x"08a0";
    tmp(01097) := x"08a0";
    tmp(01098) := x"08a0";
    tmp(01099) := x"08a0";
    tmp(01100) := x"08a0";
    tmp(01101) := x"08a0";
    tmp(01102) := x"08a0";
    tmp(01103) := x"08a0";
    tmp(01104) := x"08a0";
    tmp(01105) := x"08c0";
    tmp(01106) := x"08a0";
    tmp(01107) := x"08a0";
    tmp(01108) := x"08a0";
    tmp(01109) := x"08a0";
    tmp(01110) := x"08a0";
    tmp(01111) := x"08a0";
    tmp(01112) := x"08a0";
    tmp(01113) := x"08a0";
    tmp(01114) := x"08a0";
    tmp(01115) := x"08a0";
    tmp(01116) := x"08a0";
    tmp(01117) := x"08a0";
    tmp(01118) := x"08a0";
    tmp(01119) := x"08a0";
    tmp(01120) := x"08a0";
    tmp(01121) := x"08a0";
    tmp(01122) := x"08a0";
    tmp(01123) := x"08a0";
    tmp(01124) := x"08a0";
    tmp(01125) := x"08a0";
    tmp(01126) := x"08a0";
    tmp(01127) := x"08a0";
    tmp(01128) := x"08a0";
    tmp(01129) := x"08a0";
    tmp(01130) := x"0880";
    tmp(01131) := x"0880";
    tmp(01132) := x"0880";
    tmp(01133) := x"0880";
    tmp(01134) := x"0880";
    tmp(01135) := x"0880";
    tmp(01136) := x"0880";
    tmp(01137) := x"0880";
    tmp(01138) := x"0880";
    tmp(01139) := x"0880";
    tmp(01140) := x"0880";
    tmp(01141) := x"0880";
    tmp(01142) := x"0880";
    tmp(01143) := x"0880";
    tmp(01144) := x"0880";
    tmp(01145) := x"0880";
    tmp(01146) := x"0880";
    tmp(01147) := x"0880";
    tmp(01148) := x"0880";
    tmp(01149) := x"0880";
    tmp(01150) := x"0880";
    tmp(01151) := x"0880";
    tmp(01152) := x"0880";
    tmp(01153) := x"0880";
    tmp(01154) := x"0880";
    tmp(01155) := x"0880";
    tmp(01156) := x"0880";
    tmp(01157) := x"ffff";
    tmp(01158) := x"ffff";
    tmp(01159) := x"ffff";
    tmp(01160) := x"ffff";
    tmp(01161) := x"ffff";
    tmp(01162) := x"ffff";
    tmp(01163) := x"ffff";
    tmp(01164) := x"ffff";
    tmp(01165) := x"ffff";
    tmp(01166) := x"ffff";
    tmp(01167) := x"ffff";
    tmp(01168) := x"ffff";
    tmp(01169) := x"ffff";
    tmp(01170) := x"ffff";
    tmp(01171) := x"ffff";
    tmp(01172) := x"ffff";
    tmp(01173) := x"ffff";
    tmp(01174) := x"ffff";
    tmp(01175) := x"ffff";
    tmp(01176) := x"ffff";
    tmp(01177) := x"ffff";
    tmp(01178) := x"ffff";
    tmp(01179) := x"ffff";
    tmp(01180) := x"ffff";
    tmp(01181) := x"ffff";
    tmp(01182) := x"ffff";
    tmp(01183) := x"ffff";
    tmp(01184) := x"ffff";
    tmp(01185) := x"ffff";
    tmp(01186) := x"ffff";
    tmp(01187) := x"ffff";
    tmp(01188) := x"ffff";
    tmp(01189) := x"ffff";
    tmp(01190) := x"ffff";
    tmp(01191) := x"ffff";
    tmp(01192) := x"ffff";
    tmp(01193) := x"ffff";
    tmp(01194) := x"ffff";
    tmp(01195) := x"ffff";
    tmp(01196) := x"ffff";
    tmp(01197) := x"0820";
    tmp(01198) := x"0820";
    tmp(01199) := x"0820";
    tmp(01200) := x"0000";
    tmp(01201) := x"0020";
    tmp(01202) := x"0000";
    tmp(01203) := x"0020";
    tmp(01204) := x"0020";
    tmp(01205) := x"0020";
    tmp(01206) := x"0020";
    tmp(01207) := x"0020";
    tmp(01208) := x"0020";
    tmp(01209) := x"0020";
    tmp(01210) := x"0020";
    tmp(01211) := x"0020";
    tmp(01212) := x"0020";
    tmp(01213) := x"0020";
    tmp(01214) := x"0040";
    tmp(01215) := x"0040";
    tmp(01216) := x"0040";
    tmp(01217) := x"0040";
    tmp(01218) := x"0040";
    tmp(01219) := x"0040";
    tmp(01220) := x"0040";
    tmp(01221) := x"0040";
    tmp(01222) := x"0040";
    tmp(01223) := x"0040";
    tmp(01224) := x"0040";
    tmp(01225) := x"0040";
    tmp(01226) := x"0040";
    tmp(01227) := x"0040";
    tmp(01228) := x"0040";
    tmp(01229) := x"0040";
    tmp(01230) := x"0040";
    tmp(01231) := x"0040";
    tmp(01232) := x"0040";
    tmp(01233) := x"0040";
    tmp(01234) := x"0040";
    tmp(01235) := x"0040";
    tmp(01236) := x"0040";
    tmp(01237) := x"0040";
    tmp(01238) := x"0040";
    tmp(01239) := x"0040";
    tmp(01240) := x"0020";
    tmp(01241) := x"0040";
    tmp(01242) := x"0020";
    tmp(01243) := x"0040";
    tmp(01244) := x"0040";
    tmp(01245) := x"0040";
    tmp(01246) := x"0040";
    tmp(01247) := x"0040";
    tmp(01248) := x"0040";
    tmp(01249) := x"0040";
    tmp(01250) := x"0040";
    tmp(01251) := x"0040";
    tmp(01252) := x"0040";
    tmp(01253) := x"0040";
    tmp(01254) := x"0040";
    tmp(01255) := x"0060";
    tmp(01256) := x"0060";
    tmp(01257) := x"0060";
    tmp(01258) := x"0060";
    tmp(01259) := x"0060";
    tmp(01260) := x"0080";
    tmp(01261) := x"0880";
    tmp(01262) := x"0880";
    tmp(01263) := x"0880";
    tmp(01264) := x"08a0";
    tmp(01265) := x"08a0";
    tmp(01266) := x"08a0";
    tmp(01267) := x"08a0";
    tmp(01268) := x"08a0";
    tmp(01269) := x"08a0";
    tmp(01270) := x"0880";
    tmp(01271) := x"0880";
    tmp(01272) := x"0880";
    tmp(01273) := x"0880";
    tmp(01274) := x"0880";
    tmp(01275) := x"0880";
    tmp(01276) := x"0880";
    tmp(01277) := x"0860";
    tmp(01278) := x"0860";
    tmp(01279) := x"0860";
    tmp(01280) := x"0860";
    tmp(01281) := x"0860";
    tmp(01282) := x"0860";
    tmp(01283) := x"0860";
    tmp(01284) := x"0860";
    tmp(01285) := x"0860";
    tmp(01286) := x"0860";
    tmp(01287) := x"0860";
    tmp(01288) := x"0860";
    tmp(01289) := x"0860";
    tmp(01290) := x"0860";
    tmp(01291) := x"0860";
    tmp(01292) := x"0880";
    tmp(01293) := x"0880";
    tmp(01294) := x"0880";
    tmp(01295) := x"0880";
    tmp(01296) := x"0880";
    tmp(01297) := x"0880";
    tmp(01298) := x"0880";
    tmp(01299) := x"0880";
    tmp(01300) := x"0880";
    tmp(01301) := x"0880";
    tmp(01302) := x"0880";
    tmp(01303) := x"0060";
    tmp(01304) := x"0060";
    tmp(01305) := x"0060";
    tmp(01306) := x"0060";
    tmp(01307) := x"0060";
    tmp(01308) := x"0060";
    tmp(01309) := x"0060";
    tmp(01310) := x"0060";
    tmp(01311) := x"0080";
    tmp(01312) := x"0080";
    tmp(01313) := x"0080";
    tmp(01314) := x"0080";
    tmp(01315) := x"0080";
    tmp(01316) := x"0080";
    tmp(01317) := x"0080";
    tmp(01318) := x"0080";
    tmp(01319) := x"0080";
    tmp(01320) := x"0080";
    tmp(01321) := x"0080";
    tmp(01322) := x"0080";
    tmp(01323) := x"00a0";
    tmp(01324) := x"00a0";
    tmp(01325) := x"00a0";
    tmp(01326) := x"00a0";
    tmp(01327) := x"00a0";
    tmp(01328) := x"00a0";
    tmp(01329) := x"00a0";
    tmp(01330) := x"00a0";
    tmp(01331) := x"08a0";
    tmp(01332) := x"08a0";
    tmp(01333) := x"08a0";
    tmp(01334) := x"08a0";
    tmp(01335) := x"08a0";
    tmp(01336) := x"08a0";
    tmp(01337) := x"08a0";
    tmp(01338) := x"08a0";
    tmp(01339) := x"08a0";
    tmp(01340) := x"08a0";
    tmp(01341) := x"08a0";
    tmp(01342) := x"08c0";
    tmp(01343) := x"08c0";
    tmp(01344) := x"08a0";
    tmp(01345) := x"08c0";
    tmp(01346) := x"08a0";
    tmp(01347) := x"08c0";
    tmp(01348) := x"08a0";
    tmp(01349) := x"08a0";
    tmp(01350) := x"08c0";
    tmp(01351) := x"08c0";
    tmp(01352) := x"08a0";
    tmp(01353) := x"08a0";
    tmp(01354) := x"08a0";
    tmp(01355) := x"08a0";
    tmp(01356) := x"08a0";
    tmp(01357) := x"08a0";
    tmp(01358) := x"08a0";
    tmp(01359) := x"08a0";
    tmp(01360) := x"08a0";
    tmp(01361) := x"08a0";
    tmp(01362) := x"08a0";
    tmp(01363) := x"08a0";
    tmp(01364) := x"08a0";
    tmp(01365) := x"08a0";
    tmp(01366) := x"08a0";
    tmp(01367) := x"08a0";
    tmp(01368) := x"08a0";
    tmp(01369) := x"08a0";
    tmp(01370) := x"08a0";
    tmp(01371) := x"08a0";
    tmp(01372) := x"0880";
    tmp(01373) := x"0880";
    tmp(01374) := x"0880";
    tmp(01375) := x"0880";
    tmp(01376) := x"0880";
    tmp(01377) := x"0880";
    tmp(01378) := x"0880";
    tmp(01379) := x"0880";
    tmp(01380) := x"0880";
    tmp(01381) := x"0880";
    tmp(01382) := x"0880";
    tmp(01383) := x"0880";
    tmp(01384) := x"0880";
    tmp(01385) := x"0880";
    tmp(01386) := x"0880";
    tmp(01387) := x"0880";
    tmp(01388) := x"0880";
    tmp(01389) := x"0880";
    tmp(01390) := x"0860";
    tmp(01391) := x"0860";
    tmp(01392) := x"0860";
    tmp(01393) := x"0860";
    tmp(01394) := x"0860";
    tmp(01395) := x"0860";
    tmp(01396) := x"0860";
    tmp(01397) := x"ffff";
    tmp(01398) := x"ffff";
    tmp(01399) := x"ffff";
    tmp(01400) := x"ffff";
    tmp(01401) := x"ffff";
    tmp(01402) := x"ffff";
    tmp(01403) := x"ffff";
    tmp(01404) := x"ffff";
    tmp(01405) := x"ffff";
    tmp(01406) := x"ffff";
    tmp(01407) := x"ffff";
    tmp(01408) := x"ffff";
    tmp(01409) := x"ffff";
    tmp(01410) := x"ffff";
    tmp(01411) := x"ffff";
    tmp(01412) := x"ffff";
    tmp(01413) := x"ffff";
    tmp(01414) := x"ffff";
    tmp(01415) := x"ffff";
    tmp(01416) := x"ffff";
    tmp(01417) := x"ffff";
    tmp(01418) := x"ffff";
    tmp(01419) := x"ffff";
    tmp(01420) := x"ffff";
    tmp(01421) := x"ffff";
    tmp(01422) := x"ffff";
    tmp(01423) := x"ffff";
    tmp(01424) := x"ffff";
    tmp(01425) := x"ffff";
    tmp(01426) := x"ffff";
    tmp(01427) := x"ffff";
    tmp(01428) := x"ffff";
    tmp(01429) := x"ffff";
    tmp(01430) := x"ffff";
    tmp(01431) := x"ffff";
    tmp(01432) := x"ffff";
    tmp(01433) := x"ffff";
    tmp(01434) := x"ffff";
    tmp(01435) := x"ffff";
    tmp(01436) := x"ffff";
    tmp(01437) := x"0820";
    tmp(01438) := x"0820";
    tmp(01439) := x"0020";
    tmp(01440) := x"0000";
    tmp(01441) := x"0020";
    tmp(01442) := x"0020";
    tmp(01443) := x"0020";
    tmp(01444) := x"0020";
    tmp(01445) := x"0020";
    tmp(01446) := x"0020";
    tmp(01447) := x"0020";
    tmp(01448) := x"0020";
    tmp(01449) := x"0020";
    tmp(01450) := x"0020";
    tmp(01451) := x"0020";
    tmp(01452) := x"0020";
    tmp(01453) := x"0040";
    tmp(01454) := x"0040";
    tmp(01455) := x"0040";
    tmp(01456) := x"0040";
    tmp(01457) := x"0040";
    tmp(01458) := x"0040";
    tmp(01459) := x"0040";
    tmp(01460) := x"0040";
    tmp(01461) := x"0040";
    tmp(01462) := x"0040";
    tmp(01463) := x"0040";
    tmp(01464) := x"0040";
    tmp(01465) := x"0020";
    tmp(01466) := x"0040";
    tmp(01467) := x"0040";
    tmp(01468) := x"0040";
    tmp(01469) := x"0040";
    tmp(01470) := x"0040";
    tmp(01471) := x"0040";
    tmp(01472) := x"0040";
    tmp(01473) := x"0040";
    tmp(01474) := x"0040";
    tmp(01475) := x"0040";
    tmp(01476) := x"0040";
    tmp(01477) := x"0040";
    tmp(01478) := x"0040";
    tmp(01479) := x"0040";
    tmp(01480) := x"0040";
    tmp(01481) := x"0040";
    tmp(01482) := x"0040";
    tmp(01483) := x"0040";
    tmp(01484) := x"0040";
    tmp(01485) := x"0040";
    tmp(01486) := x"0040";
    tmp(01487) := x"0040";
    tmp(01488) := x"0040";
    tmp(01489) := x"0040";
    tmp(01490) := x"0040";
    tmp(01491) := x"0040";
    tmp(01492) := x"0040";
    tmp(01493) := x"0060";
    tmp(01494) := x"0060";
    tmp(01495) := x"0060";
    tmp(01496) := x"0060";
    tmp(01497) := x"0060";
    tmp(01498) := x"0080";
    tmp(01499) := x"0080";
    tmp(01500) := x"0880";
    tmp(01501) := x"0880";
    tmp(01502) := x"0880";
    tmp(01503) := x"0880";
    tmp(01504) := x"0880";
    tmp(01505) := x"0880";
    tmp(01506) := x"0880";
    tmp(01507) := x"0880";
    tmp(01508) := x"0880";
    tmp(01509) := x"0880";
    tmp(01510) := x"0880";
    tmp(01511) := x"0880";
    tmp(01512) := x"0880";
    tmp(01513) := x"0860";
    tmp(01514) := x"0860";
    tmp(01515) := x"0860";
    tmp(01516) := x"0860";
    tmp(01517) := x"0860";
    tmp(01518) := x"0860";
    tmp(01519) := x"0860";
    tmp(01520) := x"0860";
    tmp(01521) := x"0860";
    tmp(01522) := x"0860";
    tmp(01523) := x"0860";
    tmp(01524) := x"0860";
    tmp(01525) := x"0860";
    tmp(01526) := x"0860";
    tmp(01527) := x"0860";
    tmp(01528) := x"0860";
    tmp(01529) := x"0860";
    tmp(01530) := x"0860";
    tmp(01531) := x"0860";
    tmp(01532) := x"0880";
    tmp(01533) := x"0880";
    tmp(01534) := x"0880";
    tmp(01535) := x"0880";
    tmp(01536) := x"0880";
    tmp(01537) := x"0880";
    tmp(01538) := x"0880";
    tmp(01539) := x"0880";
    tmp(01540) := x"0880";
    tmp(01541) := x"0880";
    tmp(01542) := x"0880";
    tmp(01543) := x"0880";
    tmp(01544) := x"0060";
    tmp(01545) := x"0060";
    tmp(01546) := x"0080";
    tmp(01547) := x"0080";
    tmp(01548) := x"0060";
    tmp(01549) := x"0060";
    tmp(01550) := x"0080";
    tmp(01551) := x"0080";
    tmp(01552) := x"0080";
    tmp(01553) := x"0080";
    tmp(01554) := x"0080";
    tmp(01555) := x"0080";
    tmp(01556) := x"0080";
    tmp(01557) := x"0080";
    tmp(01558) := x"0080";
    tmp(01559) := x"0080";
    tmp(01560) := x"0080";
    tmp(01561) := x"0080";
    tmp(01562) := x"00a0";
    tmp(01563) := x"0080";
    tmp(01564) := x"00a0";
    tmp(01565) := x"00a0";
    tmp(01566) := x"00a0";
    tmp(01567) := x"00a0";
    tmp(01568) := x"00a0";
    tmp(01569) := x"00a0";
    tmp(01570) := x"00a0";
    tmp(01571) := x"00a0";
    tmp(01572) := x"00a0";
    tmp(01573) := x"00a0";
    tmp(01574) := x"08a0";
    tmp(01575) := x"08a0";
    tmp(01576) := x"08a0";
    tmp(01577) := x"08a0";
    tmp(01578) := x"08a0";
    tmp(01579) := x"08c0";
    tmp(01580) := x"08a0";
    tmp(01581) := x"08a0";
    tmp(01582) := x"08c0";
    tmp(01583) := x"08c0";
    tmp(01584) := x"08c0";
    tmp(01585) := x"08a0";
    tmp(01586) := x"08a0";
    tmp(01587) := x"08c0";
    tmp(01588) := x"08c0";
    tmp(01589) := x"08c0";
    tmp(01590) := x"08a0";
    tmp(01591) := x"08c0";
    tmp(01592) := x"08c0";
    tmp(01593) := x"08a0";
    tmp(01594) := x"08c0";
    tmp(01595) := x"08a0";
    tmp(01596) := x"08a0";
    tmp(01597) := x"08a0";
    tmp(01598) := x"08a0";
    tmp(01599) := x"08a0";
    tmp(01600) := x"08a0";
    tmp(01601) := x"08a0";
    tmp(01602) := x"08a0";
    tmp(01603) := x"08a0";
    tmp(01604) := x"08a0";
    tmp(01605) := x"08a0";
    tmp(01606) := x"08a0";
    tmp(01607) := x"08a0";
    tmp(01608) := x"08a0";
    tmp(01609) := x"08a0";
    tmp(01610) := x"08a0";
    tmp(01611) := x"08a0";
    tmp(01612) := x"08a0";
    tmp(01613) := x"0880";
    tmp(01614) := x"0880";
    tmp(01615) := x"0880";
    tmp(01616) := x"0880";
    tmp(01617) := x"0880";
    tmp(01618) := x"0880";
    tmp(01619) := x"08a0";
    tmp(01620) := x"0880";
    tmp(01621) := x"0880";
    tmp(01622) := x"0880";
    tmp(01623) := x"0880";
    tmp(01624) := x"0880";
    tmp(01625) := x"0880";
    tmp(01626) := x"0880";
    tmp(01627) := x"0880";
    tmp(01628) := x"0880";
    tmp(01629) := x"0860";
    tmp(01630) := x"0860";
    tmp(01631) := x"0860";
    tmp(01632) := x"0860";
    tmp(01633) := x"0860";
    tmp(01634) := x"0860";
    tmp(01635) := x"0860";
    tmp(01636) := x"0860";
    tmp(01637) := x"ffff";
    tmp(01638) := x"ffff";
    tmp(01639) := x"ffff";
    tmp(01640) := x"ffff";
    tmp(01641) := x"ffff";
    tmp(01642) := x"ffff";
    tmp(01643) := x"ffff";
    tmp(01644) := x"ffff";
    tmp(01645) := x"ffff";
    tmp(01646) := x"ffff";
    tmp(01647) := x"ffff";
    tmp(01648) := x"ffff";
    tmp(01649) := x"ffff";
    tmp(01650) := x"ffff";
    tmp(01651) := x"ffff";
    tmp(01652) := x"ffff";
    tmp(01653) := x"ffff";
    tmp(01654) := x"ffff";
    tmp(01655) := x"ffff";
    tmp(01656) := x"ffff";
    tmp(01657) := x"ffff";
    tmp(01658) := x"ffff";
    tmp(01659) := x"ffff";
    tmp(01660) := x"ffff";
    tmp(01661) := x"ffff";
    tmp(01662) := x"ffff";
    tmp(01663) := x"ffff";
    tmp(01664) := x"ffff";
    tmp(01665) := x"ffff";
    tmp(01666) := x"ffff";
    tmp(01667) := x"ffff";
    tmp(01668) := x"ffff";
    tmp(01669) := x"ffff";
    tmp(01670) := x"ffff";
    tmp(01671) := x"ffff";
    tmp(01672) := x"ffff";
    tmp(01673) := x"ffff";
    tmp(01674) := x"ffff";
    tmp(01675) := x"ffff";
    tmp(01676) := x"ffff";
    tmp(01677) := x"0820";
    tmp(01678) := x"0820";
    tmp(01679) := x"0020";
    tmp(01680) := x"0000";
    tmp(01681) := x"0020";
    tmp(01682) := x"0020";
    tmp(01683) := x"0020";
    tmp(01684) := x"0020";
    tmp(01685) := x"0020";
    tmp(01686) := x"0020";
    tmp(01687) := x"0020";
    tmp(01688) := x"0020";
    tmp(01689) := x"0020";
    tmp(01690) := x"0020";
    tmp(01691) := x"0020";
    tmp(01692) := x"0040";
    tmp(01693) := x"0040";
    tmp(01694) := x"0040";
    tmp(01695) := x"0040";
    tmp(01696) := x"0040";
    tmp(01697) := x"0040";
    tmp(01698) := x"0040";
    tmp(01699) := x"0040";
    tmp(01700) := x"0040";
    tmp(01701) := x"0040";
    tmp(01702) := x"0040";
    tmp(01703) := x"0040";
    tmp(01704) := x"0040";
    tmp(01705) := x"0020";
    tmp(01706) := x"0040";
    tmp(01707) := x"0040";
    tmp(01708) := x"0040";
    tmp(01709) := x"0040";
    tmp(01710) := x"0040";
    tmp(01711) := x"0040";
    tmp(01712) := x"0040";
    tmp(01713) := x"0040";
    tmp(01714) := x"0040";
    tmp(01715) := x"0040";
    tmp(01716) := x"0040";
    tmp(01717) := x"0040";
    tmp(01718) := x"0040";
    tmp(01719) := x"0040";
    tmp(01720) := x"0040";
    tmp(01721) := x"0040";
    tmp(01722) := x"0040";
    tmp(01723) := x"0040";
    tmp(01724) := x"0040";
    tmp(01725) := x"0040";
    tmp(01726) := x"0040";
    tmp(01727) := x"0040";
    tmp(01728) := x"0040";
    tmp(01729) := x"0040";
    tmp(01730) := x"0060";
    tmp(01731) := x"0060";
    tmp(01732) := x"0060";
    tmp(01733) := x"0060";
    tmp(01734) := x"0060";
    tmp(01735) := x"0060";
    tmp(01736) := x"0080";
    tmp(01737) := x"0080";
    tmp(01738) := x"0080";
    tmp(01739) := x"0880";
    tmp(01740) := x"0880";
    tmp(01741) := x"0880";
    tmp(01742) := x"0880";
    tmp(01743) := x"0880";
    tmp(01744) := x"0880";
    tmp(01745) := x"0880";
    tmp(01746) := x"0880";
    tmp(01747) := x"0880";
    tmp(01748) := x"0880";
    tmp(01749) := x"0880";
    tmp(01750) := x"0860";
    tmp(01751) := x"0880";
    tmp(01752) := x"0860";
    tmp(01753) := x"0860";
    tmp(01754) := x"0860";
    tmp(01755) := x"0860";
    tmp(01756) := x"0860";
    tmp(01757) := x"0860";
    tmp(01758) := x"0860";
    tmp(01759) := x"0860";
    tmp(01760) := x"0860";
    tmp(01761) := x"0840";
    tmp(01762) := x"0840";
    tmp(01763) := x"0840";
    tmp(01764) := x"0840";
    tmp(01765) := x"0840";
    tmp(01766) := x"0840";
    tmp(01767) := x"0840";
    tmp(01768) := x"0860";
    tmp(01769) := x"0860";
    tmp(01770) := x"0860";
    tmp(01771) := x"0860";
    tmp(01772) := x"0860";
    tmp(01773) := x"0880";
    tmp(01774) := x"0880";
    tmp(01775) := x"0880";
    tmp(01776) := x"0880";
    tmp(01777) := x"0880";
    tmp(01778) := x"0880";
    tmp(01779) := x"0880";
    tmp(01780) := x"0880";
    tmp(01781) := x"0880";
    tmp(01782) := x"0880";
    tmp(01783) := x"0880";
    tmp(01784) := x"0880";
    tmp(01785) := x"0060";
    tmp(01786) := x"0060";
    tmp(01787) := x"0880";
    tmp(01788) := x"0080";
    tmp(01789) := x"0080";
    tmp(01790) := x"0080";
    tmp(01791) := x"0080";
    tmp(01792) := x"0080";
    tmp(01793) := x"0080";
    tmp(01794) := x"0080";
    tmp(01795) := x"0080";
    tmp(01796) := x"0080";
    tmp(01797) := x"0080";
    tmp(01798) := x"0080";
    tmp(01799) := x"00a0";
    tmp(01800) := x"00a0";
    tmp(01801) := x"0080";
    tmp(01802) := x"00a0";
    tmp(01803) := x"00a0";
    tmp(01804) := x"00a0";
    tmp(01805) := x"00a0";
    tmp(01806) := x"00a0";
    tmp(01807) := x"00a0";
    tmp(01808) := x"00a0";
    tmp(01809) := x"00a0";
    tmp(01810) := x"00a0";
    tmp(01811) := x"00a0";
    tmp(01812) := x"00a0";
    tmp(01813) := x"00a0";
    tmp(01814) := x"08a0";
    tmp(01815) := x"08c0";
    tmp(01816) := x"00a0";
    tmp(01817) := x"00a0";
    tmp(01818) := x"08c0";
    tmp(01819) := x"08a0";
    tmp(01820) := x"08c0";
    tmp(01821) := x"08c0";
    tmp(01822) := x"08c0";
    tmp(01823) := x"08c0";
    tmp(01824) := x"08c0";
    tmp(01825) := x"08c0";
    tmp(01826) := x"08c0";
    tmp(01827) := x"08c0";
    tmp(01828) := x"08c0";
    tmp(01829) := x"08c0";
    tmp(01830) := x"08c0";
    tmp(01831) := x"08c0";
    tmp(01832) := x"08c0";
    tmp(01833) := x"08c0";
    tmp(01834) := x"08c0";
    tmp(01835) := x"08a0";
    tmp(01836) := x"08a0";
    tmp(01837) := x"08a0";
    tmp(01838) := x"08a0";
    tmp(01839) := x"08a0";
    tmp(01840) := x"08a0";
    tmp(01841) := x"08a0";
    tmp(01842) := x"08a0";
    tmp(01843) := x"08a0";
    tmp(01844) := x"08a0";
    tmp(01845) := x"08a0";
    tmp(01846) := x"08a0";
    tmp(01847) := x"08a0";
    tmp(01848) := x"08a0";
    tmp(01849) := x"08a0";
    tmp(01850) := x"08a0";
    tmp(01851) := x"08a0";
    tmp(01852) := x"08a0";
    tmp(01853) := x"08a0";
    tmp(01854) := x"08a0";
    tmp(01855) := x"08a0";
    tmp(01856) := x"08a0";
    tmp(01857) := x"08a0";
    tmp(01858) := x"08a0";
    tmp(01859) := x"0880";
    tmp(01860) := x"0880";
    tmp(01861) := x"0880";
    tmp(01862) := x"0880";
    tmp(01863) := x"0880";
    tmp(01864) := x"0880";
    tmp(01865) := x"0880";
    tmp(01866) := x"0880";
    tmp(01867) := x"0880";
    tmp(01868) := x"0880";
    tmp(01869) := x"0880";
    tmp(01870) := x"0860";
    tmp(01871) := x"0860";
    tmp(01872) := x"0860";
    tmp(01873) := x"0860";
    tmp(01874) := x"0860";
    tmp(01875) := x"0860";
    tmp(01876) := x"0860";
    tmp(01877) := x"ffff";
    tmp(01878) := x"ffff";
    tmp(01879) := x"ffff";
    tmp(01880) := x"ffff";
    tmp(01881) := x"ffff";
    tmp(01882) := x"ffff";
    tmp(01883) := x"ffff";
    tmp(01884) := x"ffff";
    tmp(01885) := x"ffff";
    tmp(01886) := x"ffff";
    tmp(01887) := x"ffff";
    tmp(01888) := x"ffff";
    tmp(01889) := x"ffff";
    tmp(01890) := x"ffff";
    tmp(01891) := x"ffff";
    tmp(01892) := x"ffff";
    tmp(01893) := x"ffff";
    tmp(01894) := x"ffff";
    tmp(01895) := x"ffff";
    tmp(01896) := x"ffff";
    tmp(01897) := x"ffff";
    tmp(01898) := x"ffff";
    tmp(01899) := x"ffff";
    tmp(01900) := x"ffff";
    tmp(01901) := x"ffff";
    tmp(01902) := x"ffff";
    tmp(01903) := x"ffff";
    tmp(01904) := x"ffff";
    tmp(01905) := x"ffff";
    tmp(01906) := x"ffff";
    tmp(01907) := x"ffff";
    tmp(01908) := x"ffff";
    tmp(01909) := x"ffff";
    tmp(01910) := x"ffff";
    tmp(01911) := x"ffff";
    tmp(01912) := x"ffff";
    tmp(01913) := x"ffff";
    tmp(01914) := x"ffff";
    tmp(01915) := x"ffff";
    tmp(01916) := x"ffff";
    tmp(01917) := x"0820";
    tmp(01918) := x"0020";
    tmp(01919) := x"0020";
    tmp(01920) := x"0000";
    tmp(01921) := x"0020";
    tmp(01922) := x"0020";
    tmp(01923) := x"0020";
    tmp(01924) := x"0020";
    tmp(01925) := x"0020";
    tmp(01926) := x"0020";
    tmp(01927) := x"0020";
    tmp(01928) := x"0020";
    tmp(01929) := x"0020";
    tmp(01930) := x"0020";
    tmp(01931) := x"0040";
    tmp(01932) := x"0040";
    tmp(01933) := x"0040";
    tmp(01934) := x"0040";
    tmp(01935) := x"0040";
    tmp(01936) := x"0040";
    tmp(01937) := x"0040";
    tmp(01938) := x"0040";
    tmp(01939) := x"0040";
    tmp(01940) := x"0040";
    tmp(01941) := x"0040";
    tmp(01942) := x"0040";
    tmp(01943) := x"0040";
    tmp(01944) := x"0040";
    tmp(01945) := x"0040";
    tmp(01946) := x"0040";
    tmp(01947) := x"0040";
    tmp(01948) := x"0040";
    tmp(01949) := x"0040";
    tmp(01950) := x"0040";
    tmp(01951) := x"0040";
    tmp(01952) := x"0040";
    tmp(01953) := x"0040";
    tmp(01954) := x"0040";
    tmp(01955) := x"0040";
    tmp(01956) := x"0040";
    tmp(01957) := x"0040";
    tmp(01958) := x"0040";
    tmp(01959) := x"0040";
    tmp(01960) := x"0040";
    tmp(01961) := x"0040";
    tmp(01962) := x"0040";
    tmp(01963) := x"0040";
    tmp(01964) := x"0040";
    tmp(01965) := x"0040";
    tmp(01966) := x"0040";
    tmp(01967) := x"0040";
    tmp(01968) := x"0040";
    tmp(01969) := x"0060";
    tmp(01970) := x"0060";
    tmp(01971) := x"0060";
    tmp(01972) := x"0060";
    tmp(01973) := x"0060";
    tmp(01974) := x"0060";
    tmp(01975) := x"0080";
    tmp(01976) := x"0080";
    tmp(01977) := x"0080";
    tmp(01978) := x"0080";
    tmp(01979) := x"0880";
    tmp(01980) := x"0880";
    tmp(01981) := x"0880";
    tmp(01982) := x"0880";
    tmp(01983) := x"0880";
    tmp(01984) := x"0880";
    tmp(01985) := x"0880";
    tmp(01986) := x"0880";
    tmp(01987) := x"0880";
    tmp(01988) := x"0860";
    tmp(01989) := x"0860";
    tmp(01990) := x"0860";
    tmp(01991) := x"0860";
    tmp(01992) := x"0860";
    tmp(01993) := x"0860";
    tmp(01994) := x"0860";
    tmp(01995) := x"0860";
    tmp(01996) := x"0840";
    tmp(01997) := x"0840";
    tmp(01998) := x"0840";
    tmp(01999) := x"0840";
    tmp(02000) := x"0840";
    tmp(02001) := x"0840";
    tmp(02002) := x"0840";
    tmp(02003) := x"0840";
    tmp(02004) := x"0840";
    tmp(02005) := x"0840";
    tmp(02006) := x"0840";
    tmp(02007) := x"0840";
    tmp(02008) := x"0860";
    tmp(02009) := x"0860";
    tmp(02010) := x"0860";
    tmp(02011) := x"0860";
    tmp(02012) := x"0860";
    tmp(02013) := x"0860";
    tmp(02014) := x"0880";
    tmp(02015) := x"0880";
    tmp(02016) := x"0880";
    tmp(02017) := x"0880";
    tmp(02018) := x"0880";
    tmp(02019) := x"0880";
    tmp(02020) := x"0880";
    tmp(02021) := x"0880";
    tmp(02022) := x"0880";
    tmp(02023) := x"0880";
    tmp(02024) := x"0880";
    tmp(02025) := x"0880";
    tmp(02026) := x"0880";
    tmp(02027) := x"0060";
    tmp(02028) := x"0080";
    tmp(02029) := x"0080";
    tmp(02030) := x"0080";
    tmp(02031) := x"0080";
    tmp(02032) := x"0080";
    tmp(02033) := x"0080";
    tmp(02034) := x"0080";
    tmp(02035) := x"0080";
    tmp(02036) := x"0080";
    tmp(02037) := x"0080";
    tmp(02038) := x"0080";
    tmp(02039) := x"0080";
    tmp(02040) := x"0080";
    tmp(02041) := x"00a0";
    tmp(02042) := x"00a0";
    tmp(02043) := x"00a0";
    tmp(02044) := x"00a0";
    tmp(02045) := x"00a0";
    tmp(02046) := x"00a0";
    tmp(02047) := x"00a0";
    tmp(02048) := x"00a0";
    tmp(02049) := x"00a0";
    tmp(02050) := x"00a0";
    tmp(02051) := x"00a0";
    tmp(02052) := x"00a0";
    tmp(02053) := x"00a0";
    tmp(02054) := x"00a0";
    tmp(02055) := x"00a0";
    tmp(02056) := x"00c0";
    tmp(02057) := x"00c0";
    tmp(02058) := x"08c0";
    tmp(02059) := x"08c0";
    tmp(02060) := x"00a0";
    tmp(02061) := x"08c0";
    tmp(02062) := x"08c0";
    tmp(02063) := x"08c0";
    tmp(02064) := x"08c0";
    tmp(02065) := x"08c0";
    tmp(02066) := x"08c0";
    tmp(02067) := x"08c0";
    tmp(02068) := x"08c0";
    tmp(02069) := x"08c0";
    tmp(02070) := x"08c0";
    tmp(02071) := x"08c0";
    tmp(02072) := x"08c0";
    tmp(02073) := x"08c0";
    tmp(02074) := x"08c0";
    tmp(02075) := x"08c0";
    tmp(02076) := x"08c0";
    tmp(02077) := x"08c0";
    tmp(02078) := x"08c0";
    tmp(02079) := x"08c0";
    tmp(02080) := x"08c0";
    tmp(02081) := x"08c0";
    tmp(02082) := x"08c0";
    tmp(02083) := x"08c0";
    tmp(02084) := x"08c0";
    tmp(02085) := x"08c0";
    tmp(02086) := x"08c0";
    tmp(02087) := x"08a0";
    tmp(02088) := x"08a0";
    tmp(02089) := x"08a0";
    tmp(02090) := x"08a0";
    tmp(02091) := x"08a0";
    tmp(02092) := x"08a0";
    tmp(02093) := x"08a0";
    tmp(02094) := x"08a0";
    tmp(02095) := x"08a0";
    tmp(02096) := x"08a0";
    tmp(02097) := x"08a0";
    tmp(02098) := x"0880";
    tmp(02099) := x"0880";
    tmp(02100) := x"08a0";
    tmp(02101) := x"0880";
    tmp(02102) := x"0880";
    tmp(02103) := x"0880";
    tmp(02104) := x"0880";
    tmp(02105) := x"0880";
    tmp(02106) := x"0880";
    tmp(02107) := x"0880";
    tmp(02108) := x"0880";
    tmp(02109) := x"0880";
    tmp(02110) := x"0860";
    tmp(02111) := x"0860";
    tmp(02112) := x"0860";
    tmp(02113) := x"0860";
    tmp(02114) := x"0860";
    tmp(02115) := x"0860";
    tmp(02116) := x"0860";
    tmp(02117) := x"ffff";
    tmp(02118) := x"ffff";
    tmp(02119) := x"ffff";
    tmp(02120) := x"ffff";
    tmp(02121) := x"ffff";
    tmp(02122) := x"ffff";
    tmp(02123) := x"ffff";
    tmp(02124) := x"ffff";
    tmp(02125) := x"ffff";
    tmp(02126) := x"ffff";
    tmp(02127) := x"ffff";
    tmp(02128) := x"ffff";
    tmp(02129) := x"ffff";
    tmp(02130) := x"ffff";
    tmp(02131) := x"ffff";
    tmp(02132) := x"ffff";
    tmp(02133) := x"ffff";
    tmp(02134) := x"ffff";
    tmp(02135) := x"ffff";
    tmp(02136) := x"ffff";
    tmp(02137) := x"ffff";
    tmp(02138) := x"ffff";
    tmp(02139) := x"ffff";
    tmp(02140) := x"ffff";
    tmp(02141) := x"ffff";
    tmp(02142) := x"ffff";
    tmp(02143) := x"ffff";
    tmp(02144) := x"ffff";
    tmp(02145) := x"ffff";
    tmp(02146) := x"ffff";
    tmp(02147) := x"ffff";
    tmp(02148) := x"ffff";
    tmp(02149) := x"ffff";
    tmp(02150) := x"ffff";
    tmp(02151) := x"ffff";
    tmp(02152) := x"ffff";
    tmp(02153) := x"ffff";
    tmp(02154) := x"ffff";
    tmp(02155) := x"ffff";
    tmp(02156) := x"ffff";
    tmp(02157) := x"0820";
    tmp(02158) := x"0820";
    tmp(02159) := x"0820";
    tmp(02160) := x"0000";
    tmp(02161) := x"0020";
    tmp(02162) := x"0020";
    tmp(02163) := x"0020";
    tmp(02164) := x"0020";
    tmp(02165) := x"0020";
    tmp(02166) := x"0020";
    tmp(02167) := x"0020";
    tmp(02168) := x"0020";
    tmp(02169) := x"0020";
    tmp(02170) := x"0020";
    tmp(02171) := x"0040";
    tmp(02172) := x"0040";
    tmp(02173) := x"0040";
    tmp(02174) := x"0040";
    tmp(02175) := x"0040";
    tmp(02176) := x"0040";
    tmp(02177) := x"0040";
    tmp(02178) := x"0040";
    tmp(02179) := x"0040";
    tmp(02180) := x"0040";
    tmp(02181) := x"0040";
    tmp(02182) := x"0040";
    tmp(02183) := x"0040";
    tmp(02184) := x"0040";
    tmp(02185) := x"0040";
    tmp(02186) := x"0040";
    tmp(02187) := x"0040";
    tmp(02188) := x"0040";
    tmp(02189) := x"0040";
    tmp(02190) := x"0040";
    tmp(02191) := x"0040";
    tmp(02192) := x"0040";
    tmp(02193) := x"0040";
    tmp(02194) := x"0040";
    tmp(02195) := x"0040";
    tmp(02196) := x"0040";
    tmp(02197) := x"0040";
    tmp(02198) := x"0040";
    tmp(02199) := x"0040";
    tmp(02200) := x"0040";
    tmp(02201) := x"0040";
    tmp(02202) := x"0040";
    tmp(02203) := x"0040";
    tmp(02204) := x"0040";
    tmp(02205) := x"0040";
    tmp(02206) := x"0040";
    tmp(02207) := x"0060";
    tmp(02208) := x"0060";
    tmp(02209) := x"0060";
    tmp(02210) := x"0060";
    tmp(02211) := x"0060";
    tmp(02212) := x"0060";
    tmp(02213) := x"0060";
    tmp(02214) := x"0080";
    tmp(02215) := x"0080";
    tmp(02216) := x"0080";
    tmp(02217) := x"0880";
    tmp(02218) := x"0880";
    tmp(02219) := x"0880";
    tmp(02220) := x"0880";
    tmp(02221) := x"0880";
    tmp(02222) := x"0880";
    tmp(02223) := x"0880";
    tmp(02224) := x"0880";
    tmp(02225) := x"0880";
    tmp(02226) := x"0860";
    tmp(02227) := x"0860";
    tmp(02228) := x"0860";
    tmp(02229) := x"0860";
    tmp(02230) := x"0860";
    tmp(02231) := x"0860";
    tmp(02232) := x"0860";
    tmp(02233) := x"0860";
    tmp(02234) := x"0840";
    tmp(02235) := x"0840";
    tmp(02236) := x"0840";
    tmp(02237) := x"0840";
    tmp(02238) := x"0840";
    tmp(02239) := x"0840";
    tmp(02240) := x"0840";
    tmp(02241) := x"0840";
    tmp(02242) := x"0840";
    tmp(02243) := x"0840";
    tmp(02244) := x"0840";
    tmp(02245) := x"0840";
    tmp(02246) := x"0840";
    tmp(02247) := x"0840";
    tmp(02248) := x"0860";
    tmp(02249) := x"0860";
    tmp(02250) := x"0860";
    tmp(02251) := x"0860";
    tmp(02252) := x"0860";
    tmp(02253) := x"0860";
    tmp(02254) := x"0860";
    tmp(02255) := x"0880";
    tmp(02256) := x"0880";
    tmp(02257) := x"0880";
    tmp(02258) := x"0880";
    tmp(02259) := x"0880";
    tmp(02260) := x"0880";
    tmp(02261) := x"0880";
    tmp(02262) := x"0880";
    tmp(02263) := x"0880";
    tmp(02264) := x"0880";
    tmp(02265) := x"0880";
    tmp(02266) := x"0880";
    tmp(02267) := x"0860";
    tmp(02268) := x"0060";
    tmp(02269) := x"0080";
    tmp(02270) := x"0060";
    tmp(02271) := x"0080";
    tmp(02272) := x"0080";
    tmp(02273) := x"0080";
    tmp(02274) := x"0080";
    tmp(02275) := x"0080";
    tmp(02276) := x"0080";
    tmp(02277) := x"0080";
    tmp(02278) := x"0080";
    tmp(02279) := x"0080";
    tmp(02280) := x"00a0";
    tmp(02281) := x"00a0";
    tmp(02282) := x"00a0";
    tmp(02283) := x"00a0";
    tmp(02284) := x"00a0";
    tmp(02285) := x"00a0";
    tmp(02286) := x"00a0";
    tmp(02287) := x"00a0";
    tmp(02288) := x"00a0";
    tmp(02289) := x"00a0";
    tmp(02290) := x"00a0";
    tmp(02291) := x"00a0";
    tmp(02292) := x"00a0";
    tmp(02293) := x"00c0";
    tmp(02294) := x"00a0";
    tmp(02295) := x"00a0";
    tmp(02296) := x"00a0";
    tmp(02297) := x"00a0";
    tmp(02298) := x"00c0";
    tmp(02299) := x"00c0";
    tmp(02300) := x"00c0";
    tmp(02301) := x"00c0";
    tmp(02302) := x"00c0";
    tmp(02303) := x"08c0";
    tmp(02304) := x"00c0";
    tmp(02305) := x"00c0";
    tmp(02306) := x"08c0";
    tmp(02307) := x"08c0";
    tmp(02308) := x"08c0";
    tmp(02309) := x"08c0";
    tmp(02310) := x"08c0";
    tmp(02311) := x"08c0";
    tmp(02312) := x"08c0";
    tmp(02313) := x"08c0";
    tmp(02314) := x"08c0";
    tmp(02315) := x"08c0";
    tmp(02316) := x"08c0";
    tmp(02317) := x"08c0";
    tmp(02318) := x"08c0";
    tmp(02319) := x"08c0";
    tmp(02320) := x"08c0";
    tmp(02321) := x"08c0";
    tmp(02322) := x"08c0";
    tmp(02323) := x"08c0";
    tmp(02324) := x"08c0";
    tmp(02325) := x"08c0";
    tmp(02326) := x"08c0";
    tmp(02327) := x"08c0";
    tmp(02328) := x"08c0";
    tmp(02329) := x"08c0";
    tmp(02330) := x"08c0";
    tmp(02331) := x"08a0";
    tmp(02332) := x"08a0";
    tmp(02333) := x"08a0";
    tmp(02334) := x"08a0";
    tmp(02335) := x"08a0";
    tmp(02336) := x"08a0";
    tmp(02337) := x"08a0";
    tmp(02338) := x"08a0";
    tmp(02339) := x"08a0";
    tmp(02340) := x"08a0";
    tmp(02341) := x"08a0";
    tmp(02342) := x"08a0";
    tmp(02343) := x"0880";
    tmp(02344) := x"0880";
    tmp(02345) := x"0880";
    tmp(02346) := x"0880";
    tmp(02347) := x"0880";
    tmp(02348) := x"0880";
    tmp(02349) := x"0880";
    tmp(02350) := x"0880";
    tmp(02351) := x"0860";
    tmp(02352) := x"0860";
    tmp(02353) := x"0860";
    tmp(02354) := x"0860";
    tmp(02355) := x"0860";
    tmp(02356) := x"0860";
    tmp(02357) := x"ffff";
    tmp(02358) := x"ffff";
    tmp(02359) := x"ffff";
    tmp(02360) := x"ffff";
    tmp(02361) := x"ffff";
    tmp(02362) := x"ffff";
    tmp(02363) := x"ffff";
    tmp(02364) := x"ffff";
    tmp(02365) := x"ffff";
    tmp(02366) := x"ffff";
    tmp(02367) := x"ffff";
    tmp(02368) := x"ffff";
    tmp(02369) := x"ffff";
    tmp(02370) := x"ffff";
    tmp(02371) := x"ffff";
    tmp(02372) := x"ffff";
    tmp(02373) := x"ffff";
    tmp(02374) := x"ffff";
    tmp(02375) := x"ffff";
    tmp(02376) := x"ffff";
    tmp(02377) := x"ffff";
    tmp(02378) := x"ffff";
    tmp(02379) := x"ffff";
    tmp(02380) := x"ffff";
    tmp(02381) := x"ffff";
    tmp(02382) := x"ffff";
    tmp(02383) := x"ffff";
    tmp(02384) := x"ffff";
    tmp(02385) := x"ffff";
    tmp(02386) := x"ffff";
    tmp(02387) := x"ffff";
    tmp(02388) := x"ffff";
    tmp(02389) := x"ffff";
    tmp(02390) := x"ffff";
    tmp(02391) := x"ffff";
    tmp(02392) := x"ffff";
    tmp(02393) := x"ffff";
    tmp(02394) := x"ffff";
    tmp(02395) := x"ffff";
    tmp(02396) := x"ffff";
    tmp(02397) := x"0820";
    tmp(02398) := x"0020";
    tmp(02399) := x"0020";
    tmp(02400) := x"0000";
    tmp(02401) := x"0020";
    tmp(02402) := x"0020";
    tmp(02403) := x"0020";
    tmp(02404) := x"0020";
    tmp(02405) := x"0020";
    tmp(02406) := x"0020";
    tmp(02407) := x"0020";
    tmp(02408) := x"0020";
    tmp(02409) := x"0020";
    tmp(02410) := x"0020";
    tmp(02411) := x"0040";
    tmp(02412) := x"0040";
    tmp(02413) := x"0040";
    tmp(02414) := x"0040";
    tmp(02415) := x"0040";
    tmp(02416) := x"0040";
    tmp(02417) := x"0040";
    tmp(02418) := x"0040";
    tmp(02419) := x"0020";
    tmp(02420) := x"0020";
    tmp(02421) := x"0040";
    tmp(02422) := x"0040";
    tmp(02423) := x"0040";
    tmp(02424) := x"0040";
    tmp(02425) := x"0040";
    tmp(02426) := x"0040";
    tmp(02427) := x"0040";
    tmp(02428) := x"0040";
    tmp(02429) := x"0040";
    tmp(02430) := x"0040";
    tmp(02431) := x"0040";
    tmp(02432) := x"0040";
    tmp(02433) := x"0040";
    tmp(02434) := x"0040";
    tmp(02435) := x"0040";
    tmp(02436) := x"0040";
    tmp(02437) := x"0040";
    tmp(02438) := x"0040";
    tmp(02439) := x"0040";
    tmp(02440) := x"0040";
    tmp(02441) := x"0040";
    tmp(02442) := x"0040";
    tmp(02443) := x"0040";
    tmp(02444) := x"0060";
    tmp(02445) := x"0060";
    tmp(02446) := x"0060";
    tmp(02447) := x"0060";
    tmp(02448) := x"0060";
    tmp(02449) := x"0060";
    tmp(02450) := x"0060";
    tmp(02451) := x"0060";
    tmp(02452) := x"0080";
    tmp(02453) := x"0080";
    tmp(02454) := x"0080";
    tmp(02455) := x"0080";
    tmp(02456) := x"0080";
    tmp(02457) := x"0880";
    tmp(02458) := x"0880";
    tmp(02459) := x"0880";
    tmp(02460) := x"0880";
    tmp(02461) := x"0880";
    tmp(02462) := x"0860";
    tmp(02463) := x"0860";
    tmp(02464) := x"0860";
    tmp(02465) := x"0860";
    tmp(02466) := x"0860";
    tmp(02467) := x"0860";
    tmp(02468) := x"0860";
    tmp(02469) := x"0860";
    tmp(02470) := x"0860";
    tmp(02471) := x"0840";
    tmp(02472) := x"0840";
    tmp(02473) := x"0840";
    tmp(02474) := x"0840";
    tmp(02475) := x"0840";
    tmp(02476) := x"0840";
    tmp(02477) := x"0840";
    tmp(02478) := x"0840";
    tmp(02479) := x"0840";
    tmp(02480) := x"0840";
    tmp(02481) := x"0840";
    tmp(02482) := x"0840";
    tmp(02483) := x"0840";
    tmp(02484) := x"0840";
    tmp(02485) := x"0840";
    tmp(02486) := x"0840";
    tmp(02487) := x"0860";
    tmp(02488) := x"0860";
    tmp(02489) := x"0860";
    tmp(02490) := x"0860";
    tmp(02491) := x"0860";
    tmp(02492) := x"0860";
    tmp(02493) := x"0860";
    tmp(02494) := x"0860";
    tmp(02495) := x"0880";
    tmp(02496) := x"0880";
    tmp(02497) := x"0880";
    tmp(02498) := x"0880";
    tmp(02499) := x"0880";
    tmp(02500) := x"0880";
    tmp(02501) := x"0880";
    tmp(02502) := x"0880";
    tmp(02503) := x"0880";
    tmp(02504) := x"0880";
    tmp(02505) := x"0880";
    tmp(02506) := x"0880";
    tmp(02507) := x"0860";
    tmp(02508) := x"0860";
    tmp(02509) := x"0880";
    tmp(02510) := x"0880";
    tmp(02511) := x"0880";
    tmp(02512) := x"0080";
    tmp(02513) := x"0080";
    tmp(02514) := x"0080";
    tmp(02515) := x"0080";
    tmp(02516) := x"0080";
    tmp(02517) := x"0080";
    tmp(02518) := x"0080";
    tmp(02519) := x"0080";
    tmp(02520) := x"0080";
    tmp(02521) := x"00a0";
    tmp(02522) := x"0080";
    tmp(02523) := x"00a0";
    tmp(02524) := x"00a0";
    tmp(02525) := x"00a0";
    tmp(02526) := x"00a0";
    tmp(02527) := x"00a0";
    tmp(02528) := x"00a0";
    tmp(02529) := x"00a0";
    tmp(02530) := x"00a0";
    tmp(02531) := x"00a0";
    tmp(02532) := x"00a0";
    tmp(02533) := x"00a0";
    tmp(02534) := x"00a0";
    tmp(02535) := x"00a0";
    tmp(02536) := x"00c0";
    tmp(02537) := x"00c0";
    tmp(02538) := x"00c0";
    tmp(02539) := x"00c0";
    tmp(02540) := x"00c0";
    tmp(02541) := x"00c0";
    tmp(02542) := x"00c0";
    tmp(02543) := x"00c0";
    tmp(02544) := x"00c0";
    tmp(02545) := x"00c0";
    tmp(02546) := x"00c0";
    tmp(02547) := x"08c0";
    tmp(02548) := x"08c0";
    tmp(02549) := x"08c0";
    tmp(02550) := x"00c0";
    tmp(02551) := x"08c0";
    tmp(02552) := x"08c0";
    tmp(02553) := x"08c0";
    tmp(02554) := x"08c0";
    tmp(02555) := x"08c0";
    tmp(02556) := x"08c0";
    tmp(02557) := x"08c0";
    tmp(02558) := x"08c0";
    tmp(02559) := x"08c0";
    tmp(02560) := x"08c0";
    tmp(02561) := x"08c0";
    tmp(02562) := x"08c0";
    tmp(02563) := x"08c0";
    tmp(02564) := x"08c0";
    tmp(02565) := x"08c0";
    tmp(02566) := x"08c0";
    tmp(02567) := x"08c0";
    tmp(02568) := x"08c0";
    tmp(02569) := x"08c0";
    tmp(02570) := x"08c0";
    tmp(02571) := x"08c0";
    tmp(02572) := x"08c0";
    tmp(02573) := x"08c0";
    tmp(02574) := x"08c0";
    tmp(02575) := x"08c0";
    tmp(02576) := x"08c0";
    tmp(02577) := x"08a0";
    tmp(02578) := x"08a0";
    tmp(02579) := x"08a0";
    tmp(02580) := x"08a0";
    tmp(02581) := x"08a0";
    tmp(02582) := x"08a0";
    tmp(02583) := x"08a0";
    tmp(02584) := x"08a0";
    tmp(02585) := x"08a0";
    tmp(02586) := x"08a0";
    tmp(02587) := x"08a0";
    tmp(02588) := x"0880";
    tmp(02589) := x"0880";
    tmp(02590) := x"0880";
    tmp(02591) := x"0880";
    tmp(02592) := x"0880";
    tmp(02593) := x"0880";
    tmp(02594) := x"0860";
    tmp(02595) := x"0860";
    tmp(02596) := x"0860";
    tmp(02597) := x"ffff";
    tmp(02598) := x"ffff";
    tmp(02599) := x"ffff";
    tmp(02600) := x"ffff";
    tmp(02601) := x"ffff";
    tmp(02602) := x"ffff";
    tmp(02603) := x"ffff";
    tmp(02604) := x"ffff";
    tmp(02605) := x"ffff";
    tmp(02606) := x"ffff";
    tmp(02607) := x"ffff";
    tmp(02608) := x"ffff";
    tmp(02609) := x"ffff";
    tmp(02610) := x"ffff";
    tmp(02611) := x"ffff";
    tmp(02612) := x"ffff";
    tmp(02613) := x"ffff";
    tmp(02614) := x"ffff";
    tmp(02615) := x"ffff";
    tmp(02616) := x"ffff";
    tmp(02617) := x"ffff";
    tmp(02618) := x"ffff";
    tmp(02619) := x"ffff";
    tmp(02620) := x"ffff";
    tmp(02621) := x"ffff";
    tmp(02622) := x"ffff";
    tmp(02623) := x"ffff";
    tmp(02624) := x"ffff";
    tmp(02625) := x"ffff";
    tmp(02626) := x"ffff";
    tmp(02627) := x"ffff";
    tmp(02628) := x"ffff";
    tmp(02629) := x"ffff";
    tmp(02630) := x"ffff";
    tmp(02631) := x"ffff";
    tmp(02632) := x"ffff";
    tmp(02633) := x"ffff";
    tmp(02634) := x"ffff";
    tmp(02635) := x"ffff";
    tmp(02636) := x"ffff";
    tmp(02637) := x"0820";
    tmp(02638) := x"0020";
    tmp(02639) := x"0020";
    tmp(02640) := x"0000";
    tmp(02641) := x"0020";
    tmp(02642) := x"0020";
    tmp(02643) := x"0020";
    tmp(02644) := x"0020";
    tmp(02645) := x"0020";
    tmp(02646) := x"0020";
    tmp(02647) := x"0020";
    tmp(02648) := x"0020";
    tmp(02649) := x"0020";
    tmp(02650) := x"0020";
    tmp(02651) := x"0040";
    tmp(02652) := x"0040";
    tmp(02653) := x"0040";
    tmp(02654) := x"0040";
    tmp(02655) := x"0040";
    tmp(02656) := x"0040";
    tmp(02657) := x"0040";
    tmp(02658) := x"0040";
    tmp(02659) := x"0020";
    tmp(02660) := x"0020";
    tmp(02661) := x"0040";
    tmp(02662) := x"0040";
    tmp(02663) := x"0040";
    tmp(02664) := x"0040";
    tmp(02665) := x"0040";
    tmp(02666) := x"0040";
    tmp(02667) := x"0040";
    tmp(02668) := x"0040";
    tmp(02669) := x"0040";
    tmp(02670) := x"0040";
    tmp(02671) := x"0040";
    tmp(02672) := x"0040";
    tmp(02673) := x"0040";
    tmp(02674) := x"0040";
    tmp(02675) := x"0040";
    tmp(02676) := x"0040";
    tmp(02677) := x"0040";
    tmp(02678) := x"0040";
    tmp(02679) := x"0040";
    tmp(02680) := x"0040";
    tmp(02681) := x"0040";
    tmp(02682) := x"0060";
    tmp(02683) := x"0060";
    tmp(02684) := x"0060";
    tmp(02685) := x"0060";
    tmp(02686) := x"0060";
    tmp(02687) := x"0060";
    tmp(02688) := x"0060";
    tmp(02689) := x"0060";
    tmp(02690) := x"0060";
    tmp(02691) := x"0080";
    tmp(02692) := x"0080";
    tmp(02693) := x"0080";
    tmp(02694) := x"0080";
    tmp(02695) := x"0080";
    tmp(02696) := x"0880";
    tmp(02697) := x"0880";
    tmp(02698) := x"0880";
    tmp(02699) := x"0880";
    tmp(02700) := x"0880";
    tmp(02701) := x"0860";
    tmp(02702) := x"0860";
    tmp(02703) := x"0860";
    tmp(02704) := x"0860";
    tmp(02705) := x"0860";
    tmp(02706) := x"0860";
    tmp(02707) := x"0860";
    tmp(02708) := x"0860";
    tmp(02709) := x"0840";
    tmp(02710) := x"0840";
    tmp(02711) := x"0840";
    tmp(02712) := x"0840";
    tmp(02713) := x"0840";
    tmp(02714) := x"0840";
    tmp(02715) := x"0840";
    tmp(02716) := x"0840";
    tmp(02717) := x"0840";
    tmp(02718) := x"0840";
    tmp(02719) := x"0840";
    tmp(02720) := x"0840";
    tmp(02721) := x"0840";
    tmp(02722) := x"0840";
    tmp(02723) := x"0840";
    tmp(02724) := x"0840";
    tmp(02725) := x"0840";
    tmp(02726) := x"0840";
    tmp(02727) := x"0860";
    tmp(02728) := x"0860";
    tmp(02729) := x"0860";
    tmp(02730) := x"0860";
    tmp(02731) := x"0860";
    tmp(02732) := x"0860";
    tmp(02733) := x"0860";
    tmp(02734) := x"0880";
    tmp(02735) := x"0880";
    tmp(02736) := x"0880";
    tmp(02737) := x"0880";
    tmp(02738) := x"0880";
    tmp(02739) := x"0880";
    tmp(02740) := x"0880";
    tmp(02741) := x"0880";
    tmp(02742) := x"0880";
    tmp(02743) := x"0880";
    tmp(02744) := x"0880";
    tmp(02745) := x"0880";
    tmp(02746) := x"0880";
    tmp(02747) := x"0880";
    tmp(02748) := x"0880";
    tmp(02749) := x"0880";
    tmp(02750) := x"0880";
    tmp(02751) := x"0880";
    tmp(02752) := x"0880";
    tmp(02753) := x"0080";
    tmp(02754) := x"0080";
    tmp(02755) := x"0080";
    tmp(02756) := x"0080";
    tmp(02757) := x"0080";
    tmp(02758) := x"0080";
    tmp(02759) := x"0080";
    tmp(02760) := x"0080";
    tmp(02761) := x"0080";
    tmp(02762) := x"0080";
    tmp(02763) := x"00a0";
    tmp(02764) := x"0080";
    tmp(02765) := x"00a0";
    tmp(02766) := x"00a0";
    tmp(02767) := x"00a0";
    tmp(02768) := x"00a0";
    tmp(02769) := x"00a0";
    tmp(02770) := x"00a0";
    tmp(02771) := x"00a0";
    tmp(02772) := x"00a0";
    tmp(02773) := x"00a0";
    tmp(02774) := x"00a0";
    tmp(02775) := x"00a0";
    tmp(02776) := x"00a0";
    tmp(02777) := x"00a0";
    tmp(02778) := x"00a0";
    tmp(02779) := x"00a0";
    tmp(02780) := x"00a0";
    tmp(02781) := x"00c0";
    tmp(02782) := x"00c0";
    tmp(02783) := x"00c0";
    tmp(02784) := x"00c0";
    tmp(02785) := x"00c0";
    tmp(02786) := x"08c0";
    tmp(02787) := x"08c0";
    tmp(02788) := x"00c0";
    tmp(02789) := x"08c0";
    tmp(02790) := x"08c0";
    tmp(02791) := x"08c0";
    tmp(02792) := x"08e0";
    tmp(02793) := x"08c0";
    tmp(02794) := x"08c0";
    tmp(02795) := x"08c0";
    tmp(02796) := x"08c0";
    tmp(02797) := x"08c0";
    tmp(02798) := x"08c0";
    tmp(02799) := x"08c0";
    tmp(02800) := x"08c0";
    tmp(02801) := x"08c0";
    tmp(02802) := x"08c0";
    tmp(02803) := x"08c0";
    tmp(02804) := x"08c0";
    tmp(02805) := x"08c0";
    tmp(02806) := x"08c0";
    tmp(02807) := x"08c0";
    tmp(02808) := x"08c0";
    tmp(02809) := x"08c0";
    tmp(02810) := x"08e0";
    tmp(02811) := x"08c0";
    tmp(02812) := x"08c0";
    tmp(02813) := x"08c0";
    tmp(02814) := x"08c0";
    tmp(02815) := x"08c0";
    tmp(02816) := x"08c0";
    tmp(02817) := x"08c0";
    tmp(02818) := x"08c0";
    tmp(02819) := x"08c0";
    tmp(02820) := x"08a0";
    tmp(02821) := x"08c0";
    tmp(02822) := x"08a0";
    tmp(02823) := x"08a0";
    tmp(02824) := x"08a0";
    tmp(02825) := x"08a0";
    tmp(02826) := x"08a0";
    tmp(02827) := x"08a0";
    tmp(02828) := x"08a0";
    tmp(02829) := x"08a0";
    tmp(02830) := x"0880";
    tmp(02831) := x"0880";
    tmp(02832) := x"0880";
    tmp(02833) := x"0880";
    tmp(02834) := x"0880";
    tmp(02835) := x"0860";
    tmp(02836) := x"0880";
    tmp(02837) := x"ffff";
    tmp(02838) := x"ffff";
    tmp(02839) := x"ffff";
    tmp(02840) := x"ffff";
    tmp(02841) := x"ffff";
    tmp(02842) := x"ffff";
    tmp(02843) := x"ffff";
    tmp(02844) := x"ffff";
    tmp(02845) := x"ffff";
    tmp(02846) := x"ffff";
    tmp(02847) := x"ffff";
    tmp(02848) := x"ffff";
    tmp(02849) := x"ffff";
    tmp(02850) := x"ffff";
    tmp(02851) := x"ffff";
    tmp(02852) := x"ffff";
    tmp(02853) := x"ffff";
    tmp(02854) := x"ffff";
    tmp(02855) := x"ffff";
    tmp(02856) := x"ffff";
    tmp(02857) := x"ffff";
    tmp(02858) := x"ffff";
    tmp(02859) := x"ffff";
    tmp(02860) := x"ffff";
    tmp(02861) := x"ffff";
    tmp(02862) := x"ffff";
    tmp(02863) := x"ffff";
    tmp(02864) := x"ffff";
    tmp(02865) := x"ffff";
    tmp(02866) := x"ffff";
    tmp(02867) := x"ffff";
    tmp(02868) := x"ffff";
    tmp(02869) := x"ffff";
    tmp(02870) := x"ffff";
    tmp(02871) := x"ffff";
    tmp(02872) := x"ffff";
    tmp(02873) := x"ffff";
    tmp(02874) := x"ffff";
    tmp(02875) := x"ffff";
    tmp(02876) := x"ffff";
    tmp(02877) := x"0820";
    tmp(02878) := x"0020";
    tmp(02879) := x"0820";
    tmp(02880) := x"0000";
    tmp(02881) := x"0020";
    tmp(02882) := x"0020";
    tmp(02883) := x"0020";
    tmp(02884) := x"0020";
    tmp(02885) := x"0020";
    tmp(02886) := x"0020";
    tmp(02887) := x"0020";
    tmp(02888) := x"0020";
    tmp(02889) := x"0020";
    tmp(02890) := x"0040";
    tmp(02891) := x"0040";
    tmp(02892) := x"0040";
    tmp(02893) := x"0040";
    tmp(02894) := x"0040";
    tmp(02895) := x"0040";
    tmp(02896) := x"0040";
    tmp(02897) := x"0020";
    tmp(02898) := x"0020";
    tmp(02899) := x"0020";
    tmp(02900) := x"0020";
    tmp(02901) := x"0040";
    tmp(02902) := x"0040";
    tmp(02903) := x"0840";
    tmp(02904) := x"0840";
    tmp(02905) := x"0040";
    tmp(02906) := x"0040";
    tmp(02907) := x"0040";
    tmp(02908) := x"0040";
    tmp(02909) := x"0040";
    tmp(02910) := x"0040";
    tmp(02911) := x"0040";
    tmp(02912) := x"0040";
    tmp(02913) := x"0040";
    tmp(02914) := x"0040";
    tmp(02915) := x"0060";
    tmp(02916) := x"0060";
    tmp(02917) := x"0040";
    tmp(02918) := x"0040";
    tmp(02919) := x"0060";
    tmp(02920) := x"0060";
    tmp(02921) := x"0060";
    tmp(02922) := x"0060";
    tmp(02923) := x"0060";
    tmp(02924) := x"0060";
    tmp(02925) := x"0060";
    tmp(02926) := x"0060";
    tmp(02927) := x"0060";
    tmp(02928) := x"0060";
    tmp(02929) := x"0060";
    tmp(02930) := x"0080";
    tmp(02931) := x"0080";
    tmp(02932) := x"0080";
    tmp(02933) := x"0080";
    tmp(02934) := x"0080";
    tmp(02935) := x"0080";
    tmp(02936) := x"0880";
    tmp(02937) := x"0860";
    tmp(02938) := x"0860";
    tmp(02939) := x"0860";
    tmp(02940) := x"0860";
    tmp(02941) := x"0860";
    tmp(02942) := x"0860";
    tmp(02943) := x"0860";
    tmp(02944) := x"0860";
    tmp(02945) := x"0840";
    tmp(02946) := x"0840";
    tmp(02947) := x"0840";
    tmp(02948) := x"0840";
    tmp(02949) := x"0840";
    tmp(02950) := x"0840";
    tmp(02951) := x"0840";
    tmp(02952) := x"0840";
    tmp(02953) := x"0840";
    tmp(02954) := x"0840";
    tmp(02955) := x"0840";
    tmp(02956) := x"0840";
    tmp(02957) := x"0840";
    tmp(02958) := x"0840";
    tmp(02959) := x"0840";
    tmp(02960) := x"0840";
    tmp(02961) := x"0840";
    tmp(02962) := x"0840";
    tmp(02963) := x"0840";
    tmp(02964) := x"0840";
    tmp(02965) := x"0840";
    tmp(02966) := x"0840";
    tmp(02967) := x"0840";
    tmp(02968) := x"0860";
    tmp(02969) := x"0860";
    tmp(02970) := x"0860";
    tmp(02971) := x"0860";
    tmp(02972) := x"0860";
    tmp(02973) := x"0860";
    tmp(02974) := x"0860";
    tmp(02975) := x"0860";
    tmp(02976) := x"0880";
    tmp(02977) := x"0880";
    tmp(02978) := x"0880";
    tmp(02979) := x"0880";
    tmp(02980) := x"0880";
    tmp(02981) := x"0880";
    tmp(02982) := x"0880";
    tmp(02983) := x"0880";
    tmp(02984) := x"0880";
    tmp(02985) := x"0880";
    tmp(02986) := x"0880";
    tmp(02987) := x"0880";
    tmp(02988) := x"0880";
    tmp(02989) := x"0860";
    tmp(02990) := x"0860";
    tmp(02991) := x"0880";
    tmp(02992) := x"0880";
    tmp(02993) := x"0880";
    tmp(02994) := x"0880";
    tmp(02995) := x"0880";
    tmp(02996) := x"0080";
    tmp(02997) := x"0080";
    tmp(02998) := x"0080";
    tmp(02999) := x"0080";
    tmp(03000) := x"0080";
    tmp(03001) := x"0080";
    tmp(03002) := x"0080";
    tmp(03003) := x"00a0";
    tmp(03004) := x"00a0";
    tmp(03005) := x"00a0";
    tmp(03006) := x"00a0";
    tmp(03007) := x"00a0";
    tmp(03008) := x"00a0";
    tmp(03009) := x"00a0";
    tmp(03010) := x"00a0";
    tmp(03011) := x"00a0";
    tmp(03012) := x"00a0";
    tmp(03013) := x"00a0";
    tmp(03014) := x"00a0";
    tmp(03015) := x"00a0";
    tmp(03016) := x"00a0";
    tmp(03017) := x"00a0";
    tmp(03018) := x"00a0";
    tmp(03019) := x"00a0";
    tmp(03020) := x"00a0";
    tmp(03021) := x"00a0";
    tmp(03022) := x"00c0";
    tmp(03023) := x"00c0";
    tmp(03024) := x"00c0";
    tmp(03025) := x"00c0";
    tmp(03026) := x"00c0";
    tmp(03027) := x"00c0";
    tmp(03028) := x"08c0";
    tmp(03029) := x"08c0";
    tmp(03030) := x"08c0";
    tmp(03031) := x"08c0";
    tmp(03032) := x"08c0";
    tmp(03033) := x"08c0";
    tmp(03034) := x"08c0";
    tmp(03035) := x"08c0";
    tmp(03036) := x"08c0";
    tmp(03037) := x"08c0";
    tmp(03038) := x"08c0";
    tmp(03039) := x"08e0";
    tmp(03040) := x"08c0";
    tmp(03041) := x"08e0";
    tmp(03042) := x"08c0";
    tmp(03043) := x"08c0";
    tmp(03044) := x"08c0";
    tmp(03045) := x"08c0";
    tmp(03046) := x"08c0";
    tmp(03047) := x"08c0";
    tmp(03048) := x"08c0";
    tmp(03049) := x"08e0";
    tmp(03050) := x"08c0";
    tmp(03051) := x"08c0";
    tmp(03052) := x"08c0";
    tmp(03053) := x"08c0";
    tmp(03054) := x"08c0";
    tmp(03055) := x"08c0";
    tmp(03056) := x"08c0";
    tmp(03057) := x"08c0";
    tmp(03058) := x"08c0";
    tmp(03059) := x"08c0";
    tmp(03060) := x"08c0";
    tmp(03061) := x"08c0";
    tmp(03062) := x"08c0";
    tmp(03063) := x"08c0";
    tmp(03064) := x"08c0";
    tmp(03065) := x"08a0";
    tmp(03066) := x"08a0";
    tmp(03067) := x"08a0";
    tmp(03068) := x"08a0";
    tmp(03069) := x"08a0";
    tmp(03070) := x"08a0";
    tmp(03071) := x"08a0";
    tmp(03072) := x"08a0";
    tmp(03073) := x"08a0";
    tmp(03074) := x"0880";
    tmp(03075) := x"0880";
    tmp(03076) := x"0880";
    tmp(03077) := x"ffff";
    tmp(03078) := x"ffff";
    tmp(03079) := x"ffff";
    tmp(03080) := x"ffff";
    tmp(03081) := x"ffff";
    tmp(03082) := x"ffff";
    tmp(03083) := x"ffff";
    tmp(03084) := x"ffff";
    tmp(03085) := x"ffff";
    tmp(03086) := x"ffff";
    tmp(03087) := x"ffff";
    tmp(03088) := x"ffff";
    tmp(03089) := x"ffff";
    tmp(03090) := x"ffff";
    tmp(03091) := x"ffff";
    tmp(03092) := x"ffff";
    tmp(03093) := x"ffff";
    tmp(03094) := x"ffff";
    tmp(03095) := x"ffff";
    tmp(03096) := x"ffff";
    tmp(03097) := x"ffff";
    tmp(03098) := x"ffff";
    tmp(03099) := x"ffff";
    tmp(03100) := x"ffff";
    tmp(03101) := x"ffff";
    tmp(03102) := x"ffff";
    tmp(03103) := x"ffff";
    tmp(03104) := x"ffff";
    tmp(03105) := x"ffff";
    tmp(03106) := x"ffff";
    tmp(03107) := x"ffff";
    tmp(03108) := x"ffff";
    tmp(03109) := x"ffff";
    tmp(03110) := x"ffff";
    tmp(03111) := x"ffff";
    tmp(03112) := x"ffff";
    tmp(03113) := x"ffff";
    tmp(03114) := x"ffff";
    tmp(03115) := x"ffff";
    tmp(03116) := x"ffff";
    tmp(03117) := x"0820";
    tmp(03118) := x"0020";
    tmp(03119) := x"0020";
    tmp(03120) := x"0000";
    tmp(03121) := x"0020";
    tmp(03122) := x"0020";
    tmp(03123) := x"0020";
    tmp(03124) := x"0020";
    tmp(03125) := x"0020";
    tmp(03126) := x"0020";
    tmp(03127) := x"0020";
    tmp(03128) := x"0020";
    tmp(03129) := x"0020";
    tmp(03130) := x"0040";
    tmp(03131) := x"0040";
    tmp(03132) := x"0040";
    tmp(03133) := x"0040";
    tmp(03134) := x"0040";
    tmp(03135) := x"0040";
    tmp(03136) := x"0020";
    tmp(03137) := x"0020";
    tmp(03138) := x"0020";
    tmp(03139) := x"0020";
    tmp(03140) := x"0040";
    tmp(03141) := x"0040";
    tmp(03142) := x"0040";
    tmp(03143) := x"0840";
    tmp(03144) := x"0040";
    tmp(03145) := x"0040";
    tmp(03146) := x"0040";
    tmp(03147) := x"0040";
    tmp(03148) := x"0040";
    tmp(03149) := x"0040";
    tmp(03150) := x"0040";
    tmp(03151) := x"0040";
    tmp(03152) := x"0060";
    tmp(03153) := x"0060";
    tmp(03154) := x"0060";
    tmp(03155) := x"0060";
    tmp(03156) := x"0060";
    tmp(03157) := x"0060";
    tmp(03158) := x"0060";
    tmp(03159) := x"0060";
    tmp(03160) := x"0060";
    tmp(03161) := x"0060";
    tmp(03162) := x"0060";
    tmp(03163) := x"0060";
    tmp(03164) := x"0060";
    tmp(03165) := x"0060";
    tmp(03166) := x"0060";
    tmp(03167) := x"0060";
    tmp(03168) := x"0060";
    tmp(03169) := x"0060";
    tmp(03170) := x"0060";
    tmp(03171) := x"0080";
    tmp(03172) := x"0080";
    tmp(03173) := x"0080";
    tmp(03174) := x"0060";
    tmp(03175) := x"0060";
    tmp(03176) := x"0860";
    tmp(03177) := x"0860";
    tmp(03178) := x"0860";
    tmp(03179) := x"0860";
    tmp(03180) := x"0860";
    tmp(03181) := x"0860";
    tmp(03182) := x"0860";
    tmp(03183) := x"0840";
    tmp(03184) := x"0840";
    tmp(03185) := x"0840";
    tmp(03186) := x"0840";
    tmp(03187) := x"0840";
    tmp(03188) := x"0840";
    tmp(03189) := x"0840";
    tmp(03190) := x"0840";
    tmp(03191) := x"0840";
    tmp(03192) := x"0840";
    tmp(03193) := x"0840";
    tmp(03194) := x"0840";
    tmp(03195) := x"0840";
    tmp(03196) := x"0840";
    tmp(03197) := x"0840";
    tmp(03198) := x"0840";
    tmp(03199) := x"0840";
    tmp(03200) := x"0840";
    tmp(03201) := x"0840";
    tmp(03202) := x"0840";
    tmp(03203) := x"0840";
    tmp(03204) := x"0840";
    tmp(03205) := x"0840";
    tmp(03206) := x"0840";
    tmp(03207) := x"0860";
    tmp(03208) := x"0860";
    tmp(03209) := x"0860";
    tmp(03210) := x"0860";
    tmp(03211) := x"0860";
    tmp(03212) := x"0860";
    tmp(03213) := x"0860";
    tmp(03214) := x"0860";
    tmp(03215) := x"0860";
    tmp(03216) := x"0880";
    tmp(03217) := x"0880";
    tmp(03218) := x"0880";
    tmp(03219) := x"0880";
    tmp(03220) := x"0880";
    tmp(03221) := x"0880";
    tmp(03222) := x"0880";
    tmp(03223) := x"0880";
    tmp(03224) := x"0880";
    tmp(03225) := x"0860";
    tmp(03226) := x"0860";
    tmp(03227) := x"0860";
    tmp(03228) := x"0860";
    tmp(03229) := x"0860";
    tmp(03230) := x"0860";
    tmp(03231) := x"0860";
    tmp(03232) := x"0860";
    tmp(03233) := x"0880";
    tmp(03234) := x"0880";
    tmp(03235) := x"0880";
    tmp(03236) := x"08a0";
    tmp(03237) := x"08a0";
    tmp(03238) := x"0880";
    tmp(03239) := x"0880";
    tmp(03240) := x"08a0";
    tmp(03241) := x"0880";
    tmp(03242) := x"0880";
    tmp(03243) := x"0080";
    tmp(03244) := x"0080";
    tmp(03245) := x"0080";
    tmp(03246) := x"00a0";
    tmp(03247) := x"00a0";
    tmp(03248) := x"00a0";
    tmp(03249) := x"00a0";
    tmp(03250) := x"00a0";
    tmp(03251) := x"00a0";
    tmp(03252) := x"00a0";
    tmp(03253) := x"00a0";
    tmp(03254) := x"00a0";
    tmp(03255) := x"00a0";
    tmp(03256) := x"00a0";
    tmp(03257) := x"00a0";
    tmp(03258) := x"00a0";
    tmp(03259) := x"00a0";
    tmp(03260) := x"00a0";
    tmp(03261) := x"00a0";
    tmp(03262) := x"00a0";
    tmp(03263) := x"00c0";
    tmp(03264) := x"00a0";
    tmp(03265) := x"00c0";
    tmp(03266) := x"08c0";
    tmp(03267) := x"08c0";
    tmp(03268) := x"00c0";
    tmp(03269) := x"08c0";
    tmp(03270) := x"00c0";
    tmp(03271) := x"08c0";
    tmp(03272) := x"08c0";
    tmp(03273) := x"08c0";
    tmp(03274) := x"08c0";
    tmp(03275) := x"08c0";
    tmp(03276) := x"08c0";
    tmp(03277) := x"08c0";
    tmp(03278) := x"08c0";
    tmp(03279) := x"08c0";
    tmp(03280) := x"08c0";
    tmp(03281) := x"08c0";
    tmp(03282) := x"08c0";
    tmp(03283) := x"08c0";
    tmp(03284) := x"08c0";
    tmp(03285) := x"08c0";
    tmp(03286) := x"08c0";
    tmp(03287) := x"08c0";
    tmp(03288) := x"08c0";
    tmp(03289) := x"08c0";
    tmp(03290) := x"08c0";
    tmp(03291) := x"08c0";
    tmp(03292) := x"08c0";
    tmp(03293) := x"08c0";
    tmp(03294) := x"08c0";
    tmp(03295) := x"08c0";
    tmp(03296) := x"08c0";
    tmp(03297) := x"08c0";
    tmp(03298) := x"08c0";
    tmp(03299) := x"08c0";
    tmp(03300) := x"08c0";
    tmp(03301) := x"08c0";
    tmp(03302) := x"08c0";
    tmp(03303) := x"08c0";
    tmp(03304) := x"08c0";
    tmp(03305) := x"08c0";
    tmp(03306) := x"08c0";
    tmp(03307) := x"08c0";
    tmp(03308) := x"08a0";
    tmp(03309) := x"08a0";
    tmp(03310) := x"08a0";
    tmp(03311) := x"08a0";
    tmp(03312) := x"08a0";
    tmp(03313) := x"08a0";
    tmp(03314) := x"08a0";
    tmp(03315) := x"08a0";
    tmp(03316) := x"08a0";
    tmp(03317) := x"ffff";
    tmp(03318) := x"ffff";
    tmp(03319) := x"ffff";
    tmp(03320) := x"ffff";
    tmp(03321) := x"ffff";
    tmp(03322) := x"ffff";
    tmp(03323) := x"ffff";
    tmp(03324) := x"ffff";
    tmp(03325) := x"ffff";
    tmp(03326) := x"ffff";
    tmp(03327) := x"ffff";
    tmp(03328) := x"ffff";
    tmp(03329) := x"ffff";
    tmp(03330) := x"ffff";
    tmp(03331) := x"ffff";
    tmp(03332) := x"ffff";
    tmp(03333) := x"ffff";
    tmp(03334) := x"ffff";
    tmp(03335) := x"ffff";
    tmp(03336) := x"ffff";
    tmp(03337) := x"ffff";
    tmp(03338) := x"ffff";
    tmp(03339) := x"ffff";
    tmp(03340) := x"ffff";
    tmp(03341) := x"ffff";
    tmp(03342) := x"ffff";
    tmp(03343) := x"ffff";
    tmp(03344) := x"ffff";
    tmp(03345) := x"ffff";
    tmp(03346) := x"ffff";
    tmp(03347) := x"ffff";
    tmp(03348) := x"ffff";
    tmp(03349) := x"ffff";
    tmp(03350) := x"ffff";
    tmp(03351) := x"ffff";
    tmp(03352) := x"ffff";
    tmp(03353) := x"ffff";
    tmp(03354) := x"ffff";
    tmp(03355) := x"ffff";
    tmp(03356) := x"ffff";
    tmp(03357) := x"0020";
    tmp(03358) := x"0020";
    tmp(03359) := x"0020";
    tmp(03360) := x"0000";
    tmp(03361) := x"0020";
    tmp(03362) := x"0020";
    tmp(03363) := x"0020";
    tmp(03364) := x"0020";
    tmp(03365) := x"0020";
    tmp(03366) := x"0020";
    tmp(03367) := x"0020";
    tmp(03368) := x"0020";
    tmp(03369) := x"0020";
    tmp(03370) := x"0020";
    tmp(03371) := x"0040";
    tmp(03372) := x"0040";
    tmp(03373) := x"0040";
    tmp(03374) := x"0040";
    tmp(03375) := x"0020";
    tmp(03376) := x"0020";
    tmp(03377) := x"0020";
    tmp(03378) := x"0020";
    tmp(03379) := x"0040";
    tmp(03380) := x"0020";
    tmp(03381) := x"0040";
    tmp(03382) := x"0040";
    tmp(03383) := x"0840";
    tmp(03384) := x"0040";
    tmp(03385) := x"0840";
    tmp(03386) := x"0040";
    tmp(03387) := x"0040";
    tmp(03388) := x"0040";
    tmp(03389) := x"0040";
    tmp(03390) := x"0040";
    tmp(03391) := x"0060";
    tmp(03392) := x"0060";
    tmp(03393) := x"0060";
    tmp(03394) := x"0060";
    tmp(03395) := x"0060";
    tmp(03396) := x"0060";
    tmp(03397) := x"0060";
    tmp(03398) := x"0060";
    tmp(03399) := x"0060";
    tmp(03400) := x"0060";
    tmp(03401) := x"0060";
    tmp(03402) := x"0060";
    tmp(03403) := x"0060";
    tmp(03404) := x"0060";
    tmp(03405) := x"0060";
    tmp(03406) := x"0060";
    tmp(03407) := x"0060";
    tmp(03408) := x"0060";
    tmp(03409) := x"0060";
    tmp(03410) := x"0060";
    tmp(03411) := x"0060";
    tmp(03412) := x"0060";
    tmp(03413) := x"0060";
    tmp(03414) := x"0060";
    tmp(03415) := x"0860";
    tmp(03416) := x"0860";
    tmp(03417) := x"0860";
    tmp(03418) := x"0860";
    tmp(03419) := x"0860";
    tmp(03420) := x"0860";
    tmp(03421) := x"0840";
    tmp(03422) := x"0840";
    tmp(03423) := x"0840";
    tmp(03424) := x"0840";
    tmp(03425) := x"0840";
    tmp(03426) := x"0840";
    tmp(03427) := x"0840";
    tmp(03428) := x"0840";
    tmp(03429) := x"0840";
    tmp(03430) := x"0840";
    tmp(03431) := x"0840";
    tmp(03432) := x"0840";
    tmp(03433) := x"0840";
    tmp(03434) := x"0840";
    tmp(03435) := x"0840";
    tmp(03436) := x"0840";
    tmp(03437) := x"0840";
    tmp(03438) := x"0840";
    tmp(03439) := x"0840";
    tmp(03440) := x"0840";
    tmp(03441) := x"0840";
    tmp(03442) := x"0840";
    tmp(03443) := x"0840";
    tmp(03444) := x"0840";
    tmp(03445) := x"0840";
    tmp(03446) := x"0840";
    tmp(03447) := x"0860";
    tmp(03448) := x"0860";
    tmp(03449) := x"0860";
    tmp(03450) := x"0860";
    tmp(03451) := x"0860";
    tmp(03452) := x"0860";
    tmp(03453) := x"0860";
    tmp(03454) := x"0880";
    tmp(03455) := x"0880";
    tmp(03456) := x"0880";
    tmp(03457) := x"0880";
    tmp(03458) := x"0880";
    tmp(03459) := x"0880";
    tmp(03460) := x"0880";
    tmp(03461) := x"0880";
    tmp(03462) := x"0880";
    tmp(03463) := x"0860";
    tmp(03464) := x"0840";
    tmp(03465) := x"0020";
    tmp(03466) := x"0020";
    tmp(03467) := x"0020";
    tmp(03468) := x"0020";
    tmp(03469) := x"0020";
    tmp(03470) := x"0020";
    tmp(03471) := x"0020";
    tmp(03472) := x"0020";
    tmp(03473) := x"0820";
    tmp(03474) := x"0821";
    tmp(03475) := x"0841";
    tmp(03476) := x"0841";
    tmp(03477) := x"0861";
    tmp(03478) := x"0881";
    tmp(03479) := x"10a1";
    tmp(03480) := x"1922";
    tmp(03481) := x"1102";
    tmp(03482) := x"10e1";
    tmp(03483) := x"08c0";
    tmp(03484) := x"08a0";
    tmp(03485) := x"08a0";
    tmp(03486) := x"0080";
    tmp(03487) := x"0080";
    tmp(03488) := x"00a0";
    tmp(03489) := x"00a0";
    tmp(03490) := x"00a0";
    tmp(03491) := x"00a0";
    tmp(03492) := x"00a0";
    tmp(03493) := x"00a0";
    tmp(03494) := x"00a0";
    tmp(03495) := x"00a0";
    tmp(03496) := x"00a0";
    tmp(03497) := x"00a0";
    tmp(03498) := x"00a0";
    tmp(03499) := x"00a0";
    tmp(03500) := x"00a0";
    tmp(03501) := x"00a0";
    tmp(03502) := x"00a0";
    tmp(03503) := x"00a0";
    tmp(03504) := x"00a0";
    tmp(03505) := x"00a0";
    tmp(03506) := x"00c0";
    tmp(03507) := x"00c0";
    tmp(03508) := x"00c0";
    tmp(03509) := x"08c0";
    tmp(03510) := x"08c0";
    tmp(03511) := x"08c0";
    tmp(03512) := x"08c0";
    tmp(03513) := x"08c0";
    tmp(03514) := x"08c0";
    tmp(03515) := x"08c0";
    tmp(03516) := x"08c0";
    tmp(03517) := x"08c0";
    tmp(03518) := x"08c0";
    tmp(03519) := x"08c0";
    tmp(03520) := x"08c0";
    tmp(03521) := x"08c0";
    tmp(03522) := x"08c0";
    tmp(03523) := x"08c0";
    tmp(03524) := x"08e0";
    tmp(03525) := x"08c0";
    tmp(03526) := x"08c0";
    tmp(03527) := x"08c0";
    tmp(03528) := x"08c0";
    tmp(03529) := x"08c0";
    tmp(03530) := x"08c0";
    tmp(03531) := x"08c0";
    tmp(03532) := x"08c0";
    tmp(03533) := x"08c0";
    tmp(03534) := x"08c0";
    tmp(03535) := x"08c0";
    tmp(03536) := x"08c0";
    tmp(03537) := x"08c0";
    tmp(03538) := x"08c0";
    tmp(03539) := x"08c0";
    tmp(03540) := x"08c0";
    tmp(03541) := x"08c0";
    tmp(03542) := x"08c0";
    tmp(03543) := x"08c0";
    tmp(03544) := x"08c0";
    tmp(03545) := x"08c0";
    tmp(03546) := x"08c0";
    tmp(03547) := x"08c0";
    tmp(03548) := x"08a0";
    tmp(03549) := x"08c0";
    tmp(03550) := x"08a0";
    tmp(03551) := x"08a0";
    tmp(03552) := x"08a0";
    tmp(03553) := x"08a0";
    tmp(03554) := x"08a0";
    tmp(03555) := x"08a0";
    tmp(03556) := x"08a0";
    tmp(03557) := x"ffff";
    tmp(03558) := x"ffff";
    tmp(03559) := x"ffff";
    tmp(03560) := x"ffff";
    tmp(03561) := x"ffff";
    tmp(03562) := x"ffff";
    tmp(03563) := x"ffff";
    tmp(03564) := x"ffff";
    tmp(03565) := x"ffff";
    tmp(03566) := x"ffff";
    tmp(03567) := x"ffff";
    tmp(03568) := x"ffff";
    tmp(03569) := x"ffff";
    tmp(03570) := x"ffff";
    tmp(03571) := x"ffff";
    tmp(03572) := x"ffff";
    tmp(03573) := x"ffff";
    tmp(03574) := x"ffff";
    tmp(03575) := x"ffff";
    tmp(03576) := x"ffff";
    tmp(03577) := x"ffff";
    tmp(03578) := x"ffff";
    tmp(03579) := x"ffff";
    tmp(03580) := x"ffff";
    tmp(03581) := x"ffff";
    tmp(03582) := x"ffff";
    tmp(03583) := x"ffff";
    tmp(03584) := x"ffff";
    tmp(03585) := x"ffff";
    tmp(03586) := x"ffff";
    tmp(03587) := x"ffff";
    tmp(03588) := x"ffff";
    tmp(03589) := x"ffff";
    tmp(03590) := x"ffff";
    tmp(03591) := x"ffff";
    tmp(03592) := x"ffff";
    tmp(03593) := x"ffff";
    tmp(03594) := x"ffff";
    tmp(03595) := x"ffff";
    tmp(03596) := x"ffff";
    tmp(03597) := x"0020";
    tmp(03598) := x"0020";
    tmp(03599) := x"0020";
    tmp(03600) := x"0000";
    tmp(03601) := x"0020";
    tmp(03602) := x"0020";
    tmp(03603) := x"0020";
    tmp(03604) := x"0020";
    tmp(03605) := x"0020";
    tmp(03606) := x"0020";
    tmp(03607) := x"0020";
    tmp(03608) := x"0020";
    tmp(03609) := x"0020";
    tmp(03610) := x"0020";
    tmp(03611) := x"0040";
    tmp(03612) := x"0040";
    tmp(03613) := x"0040";
    tmp(03614) := x"0020";
    tmp(03615) := x"0020";
    tmp(03616) := x"0020";
    tmp(03617) := x"0020";
    tmp(03618) := x"0040";
    tmp(03619) := x"0040";
    tmp(03620) := x"0040";
    tmp(03621) := x"0040";
    tmp(03622) := x"0840";
    tmp(03623) := x"0840";
    tmp(03624) := x"0840";
    tmp(03625) := x"0840";
    tmp(03626) := x"0040";
    tmp(03627) := x"0040";
    tmp(03628) := x"0040";
    tmp(03629) := x"0040";
    tmp(03630) := x"0040";
    tmp(03631) := x"0060";
    tmp(03632) := x"0060";
    tmp(03633) := x"0060";
    tmp(03634) := x"0060";
    tmp(03635) := x"0060";
    tmp(03636) := x"0060";
    tmp(03637) := x"0060";
    tmp(03638) := x"0060";
    tmp(03639) := x"0060";
    tmp(03640) := x"0060";
    tmp(03641) := x"0060";
    tmp(03642) := x"0060";
    tmp(03643) := x"0060";
    tmp(03644) := x"0060";
    tmp(03645) := x"0060";
    tmp(03646) := x"0060";
    tmp(03647) := x"0060";
    tmp(03648) := x"0060";
    tmp(03649) := x"0060";
    tmp(03650) := x"0060";
    tmp(03651) := x"0060";
    tmp(03652) := x"0060";
    tmp(03653) := x"0860";
    tmp(03654) := x"0860";
    tmp(03655) := x"0860";
    tmp(03656) := x"0860";
    tmp(03657) := x"0860";
    tmp(03658) := x"0860";
    tmp(03659) := x"0860";
    tmp(03660) := x"0840";
    tmp(03661) := x"0840";
    tmp(03662) := x"0840";
    tmp(03663) := x"0840";
    tmp(03664) := x"0840";
    tmp(03665) := x"0840";
    tmp(03666) := x"0840";
    tmp(03667) := x"0840";
    tmp(03668) := x"0840";
    tmp(03669) := x"0840";
    tmp(03670) := x"0840";
    tmp(03671) := x"0840";
    tmp(03672) := x"0840";
    tmp(03673) := x"0840";
    tmp(03674) := x"0840";
    tmp(03675) := x"0840";
    tmp(03676) := x"0840";
    tmp(03677) := x"0840";
    tmp(03678) := x"0840";
    tmp(03679) := x"0840";
    tmp(03680) := x"0840";
    tmp(03681) := x"0840";
    tmp(03682) := x"0840";
    tmp(03683) := x"0840";
    tmp(03684) := x"0840";
    tmp(03685) := x"0840";
    tmp(03686) := x"0840";
    tmp(03687) := x"0840";
    tmp(03688) := x"0840";
    tmp(03689) := x"0860";
    tmp(03690) := x"0860";
    tmp(03691) := x"0860";
    tmp(03692) := x"0860";
    tmp(03693) := x"0860";
    tmp(03694) := x"0860";
    tmp(03695) := x"0880";
    tmp(03696) := x"0880";
    tmp(03697) := x"0880";
    tmp(03698) := x"0880";
    tmp(03699) := x"0880";
    tmp(03700) := x"0880";
    tmp(03701) := x"0880";
    tmp(03702) := x"0880";
    tmp(03703) := x"0840";
    tmp(03704) := x"0000";
    tmp(03705) := x"0000";
    tmp(03706) := x"0000";
    tmp(03707) := x"0000";
    tmp(03708) := x"0000";
    tmp(03709) := x"0000";
    tmp(03710) := x"0000";
    tmp(03711) := x"0000";
    tmp(03712) := x"0000";
    tmp(03713) := x"0000";
    tmp(03714) := x"0000";
    tmp(03715) := x"0000";
    tmp(03716) := x"0000";
    tmp(03717) := x"0020";
    tmp(03718) := x"0020";
    tmp(03719) := x"0821";
    tmp(03720) := x"0862";
    tmp(03721) := x"10a2";
    tmp(03722) := x"1903";
    tmp(03723) := x"1923";
    tmp(03724) := x"1922";
    tmp(03725) := x"1121";
    tmp(03726) := x"08e1";
    tmp(03727) := x"08a0";
    tmp(03728) := x"08a0";
    tmp(03729) := x"0080";
    tmp(03730) := x"00a0";
    tmp(03731) := x"00a0";
    tmp(03732) := x"00a0";
    tmp(03733) := x"00a0";
    tmp(03734) := x"00a0";
    tmp(03735) := x"00a0";
    tmp(03736) := x"00a0";
    tmp(03737) := x"00a0";
    tmp(03738) := x"00a0";
    tmp(03739) := x"00a0";
    tmp(03740) := x"00a0";
    tmp(03741) := x"00a0";
    tmp(03742) := x"00a0";
    tmp(03743) := x"00a0";
    tmp(03744) := x"00c0";
    tmp(03745) := x"00a0";
    tmp(03746) := x"00a0";
    tmp(03747) := x"00c0";
    tmp(03748) := x"08c0";
    tmp(03749) := x"08c0";
    tmp(03750) := x"08c0";
    tmp(03751) := x"08c0";
    tmp(03752) := x"08c0";
    tmp(03753) := x"08c0";
    tmp(03754) := x"08c0";
    tmp(03755) := x"08c0";
    tmp(03756) := x"08c0";
    tmp(03757) := x"08c0";
    tmp(03758) := x"08c0";
    tmp(03759) := x"08c0";
    tmp(03760) := x"08c0";
    tmp(03761) := x"08c0";
    tmp(03762) := x"08c0";
    tmp(03763) := x"08c0";
    tmp(03764) := x"08c0";
    tmp(03765) := x"08c0";
    tmp(03766) := x"08c0";
    tmp(03767) := x"08c0";
    tmp(03768) := x"08c0";
    tmp(03769) := x"08c0";
    tmp(03770) := x"08c0";
    tmp(03771) := x"08c0";
    tmp(03772) := x"08c0";
    tmp(03773) := x"08c0";
    tmp(03774) := x"08c0";
    tmp(03775) := x"08c0";
    tmp(03776) := x"08c0";
    tmp(03777) := x"08c0";
    tmp(03778) := x"08c0";
    tmp(03779) := x"08c0";
    tmp(03780) := x"08c0";
    tmp(03781) := x"08c0";
    tmp(03782) := x"08c0";
    tmp(03783) := x"08c0";
    tmp(03784) := x"08c0";
    tmp(03785) := x"08c0";
    tmp(03786) := x"08c0";
    tmp(03787) := x"08c0";
    tmp(03788) := x"08c0";
    tmp(03789) := x"08c0";
    tmp(03790) := x"08c0";
    tmp(03791) := x"08a0";
    tmp(03792) := x"08a0";
    tmp(03793) := x"08a0";
    tmp(03794) := x"08a0";
    tmp(03795) := x"08a0";
    tmp(03796) := x"08a0";
    tmp(03797) := x"ffff";
    tmp(03798) := x"ffff";
    tmp(03799) := x"ffff";
    tmp(03800) := x"ffff";
    tmp(03801) := x"ffff";
    tmp(03802) := x"ffff";
    tmp(03803) := x"ffff";
    tmp(03804) := x"ffff";
    tmp(03805) := x"ffff";
    tmp(03806) := x"ffff";
    tmp(03807) := x"ffff";
    tmp(03808) := x"ffff";
    tmp(03809) := x"ffff";
    tmp(03810) := x"ffff";
    tmp(03811) := x"ffff";
    tmp(03812) := x"ffff";
    tmp(03813) := x"ffff";
    tmp(03814) := x"ffff";
    tmp(03815) := x"ffff";
    tmp(03816) := x"ffff";
    tmp(03817) := x"ffff";
    tmp(03818) := x"ffff";
    tmp(03819) := x"ffff";
    tmp(03820) := x"ffff";
    tmp(03821) := x"ffff";
    tmp(03822) := x"ffff";
    tmp(03823) := x"ffff";
    tmp(03824) := x"ffff";
    tmp(03825) := x"ffff";
    tmp(03826) := x"ffff";
    tmp(03827) := x"ffff";
    tmp(03828) := x"ffff";
    tmp(03829) := x"ffff";
    tmp(03830) := x"ffff";
    tmp(03831) := x"ffff";
    tmp(03832) := x"ffff";
    tmp(03833) := x"ffff";
    tmp(03834) := x"ffff";
    tmp(03835) := x"ffff";
    tmp(03836) := x"ffff";
    tmp(03837) := x"0820";
    tmp(03838) := x"0020";
    tmp(03839) := x"0020";
    tmp(03840) := x"0000";
    tmp(03841) := x"0020";
    tmp(03842) := x"0020";
    tmp(03843) := x"0020";
    tmp(03844) := x"0020";
    tmp(03845) := x"0020";
    tmp(03846) := x"0020";
    tmp(03847) := x"0020";
    tmp(03848) := x"0020";
    tmp(03849) := x"0020";
    tmp(03850) := x"0020";
    tmp(03851) := x"0020";
    tmp(03852) := x"0040";
    tmp(03853) := x"0040";
    tmp(03854) := x"0040";
    tmp(03855) := x"0040";
    tmp(03856) := x"0020";
    tmp(03857) := x"0040";
    tmp(03858) := x"0040";
    tmp(03859) := x"0040";
    tmp(03860) := x"0040";
    tmp(03861) := x"0040";
    tmp(03862) := x"0040";
    tmp(03863) := x"0840";
    tmp(03864) := x"0840";
    tmp(03865) := x"0840";
    tmp(03866) := x"0040";
    tmp(03867) := x"0040";
    tmp(03868) := x"0040";
    tmp(03869) := x"0040";
    tmp(03870) := x"0040";
    tmp(03871) := x"0040";
    tmp(03872) := x"0060";
    tmp(03873) := x"0060";
    tmp(03874) := x"0060";
    tmp(03875) := x"0060";
    tmp(03876) := x"0060";
    tmp(03877) := x"0060";
    tmp(03878) := x"0060";
    tmp(03879) := x"0060";
    tmp(03880) := x"0060";
    tmp(03881) := x"0060";
    tmp(03882) := x"0060";
    tmp(03883) := x"0060";
    tmp(03884) := x"0060";
    tmp(03885) := x"0060";
    tmp(03886) := x"0060";
    tmp(03887) := x"0060";
    tmp(03888) := x"0060";
    tmp(03889) := x"0060";
    tmp(03890) := x"0060";
    tmp(03891) := x"0060";
    tmp(03892) := x"0860";
    tmp(03893) := x"0860";
    tmp(03894) := x"0860";
    tmp(03895) := x"0860";
    tmp(03896) := x"0860";
    tmp(03897) := x"0860";
    tmp(03898) := x"0840";
    tmp(03899) := x"0840";
    tmp(03900) := x"0840";
    tmp(03901) := x"0840";
    tmp(03902) := x"0840";
    tmp(03903) := x"0840";
    tmp(03904) := x"0840";
    tmp(03905) := x"0840";
    tmp(03906) := x"0840";
    tmp(03907) := x"0820";
    tmp(03908) := x"0840";
    tmp(03909) := x"0840";
    tmp(03910) := x"0840";
    tmp(03911) := x"0840";
    tmp(03912) := x"0840";
    tmp(03913) := x"0840";
    tmp(03914) := x"0840";
    tmp(03915) := x"0840";
    tmp(03916) := x"0840";
    tmp(03917) := x"0840";
    tmp(03918) := x"0840";
    tmp(03919) := x"0840";
    tmp(03920) := x"0840";
    tmp(03921) := x"0840";
    tmp(03922) := x"0840";
    tmp(03923) := x"0840";
    tmp(03924) := x"0840";
    tmp(03925) := x"0840";
    tmp(03926) := x"0840";
    tmp(03927) := x"0840";
    tmp(03928) := x"0840";
    tmp(03929) := x"0860";
    tmp(03930) := x"0860";
    tmp(03931) := x"0860";
    tmp(03932) := x"0860";
    tmp(03933) := x"0860";
    tmp(03934) := x"0860";
    tmp(03935) := x"0880";
    tmp(03936) := x"0880";
    tmp(03937) := x"0880";
    tmp(03938) := x"0880";
    tmp(03939) := x"0880";
    tmp(03940) := x"0880";
    tmp(03941) := x"0880";
    tmp(03942) := x"0880";
    tmp(03943) := x"0860";
    tmp(03944) := x"0020";
    tmp(03945) := x"0020";
    tmp(03946) := x"0000";
    tmp(03947) := x"0000";
    tmp(03948) := x"0000";
    tmp(03949) := x"0000";
    tmp(03950) := x"0000";
    tmp(03951) := x"0000";
    tmp(03952) := x"0000";
    tmp(03953) := x"0000";
    tmp(03954) := x"0000";
    tmp(03955) := x"0000";
    tmp(03956) := x"0000";
    tmp(03957) := x"0000";
    tmp(03958) := x"0000";
    tmp(03959) := x"0000";
    tmp(03960) := x"0020";
    tmp(03961) := x"0821";
    tmp(03962) := x"0841";
    tmp(03963) := x"0882";
    tmp(03964) := x"10a2";
    tmp(03965) := x"18e3";
    tmp(03966) := x"1943";
    tmp(03967) := x"1922";
    tmp(03968) := x"1101";
    tmp(03969) := x"08e0";
    tmp(03970) := x"08a0";
    tmp(03971) := x"00a0";
    tmp(03972) := x"00a0";
    tmp(03973) := x"00a0";
    tmp(03974) := x"00a0";
    tmp(03975) := x"00a0";
    tmp(03976) := x"00a0";
    tmp(03977) := x"00a0";
    tmp(03978) := x"00a0";
    tmp(03979) := x"00a0";
    tmp(03980) := x"00a0";
    tmp(03981) := x"00a0";
    tmp(03982) := x"00a0";
    tmp(03983) := x"00c0";
    tmp(03984) := x"00a0";
    tmp(03985) := x"00a0";
    tmp(03986) := x"08c0";
    tmp(03987) := x"08c0";
    tmp(03988) := x"08c0";
    tmp(03989) := x"08c0";
    tmp(03990) := x"08c0";
    tmp(03991) := x"08c0";
    tmp(03992) := x"08c0";
    tmp(03993) := x"08c0";
    tmp(03994) := x"08c0";
    tmp(03995) := x"08c0";
    tmp(03996) := x"08c0";
    tmp(03997) := x"08c0";
    tmp(03998) := x"08c0";
    tmp(03999) := x"08c0";
    tmp(04000) := x"08c0";
    tmp(04001) := x"08c0";
    tmp(04002) := x"08c0";
    tmp(04003) := x"08c0";
    tmp(04004) := x"08c0";
    tmp(04005) := x"08c0";
    tmp(04006) := x"08c0";
    tmp(04007) := x"08c0";
    tmp(04008) := x"08c0";
    tmp(04009) := x"08c0";
    tmp(04010) := x"08c0";
    tmp(04011) := x"08c0";
    tmp(04012) := x"08c0";
    tmp(04013) := x"08c0";
    tmp(04014) := x"08c0";
    tmp(04015) := x"08c0";
    tmp(04016) := x"08c0";
    tmp(04017) := x"08c0";
    tmp(04018) := x"08c0";
    tmp(04019) := x"08c0";
    tmp(04020) := x"08c0";
    tmp(04021) := x"08c0";
    tmp(04022) := x"08c0";
    tmp(04023) := x"08c0";
    tmp(04024) := x"08c0";
    tmp(04025) := x"08c0";
    tmp(04026) := x"08c0";
    tmp(04027) := x"08c0";
    tmp(04028) := x"08a0";
    tmp(04029) := x"08a0";
    tmp(04030) := x"08a0";
    tmp(04031) := x"08a0";
    tmp(04032) := x"08a0";
    tmp(04033) := x"08a0";
    tmp(04034) := x"08a0";
    tmp(04035) := x"08a0";
    tmp(04036) := x"08a0";
    tmp(04037) := x"ffff";
    tmp(04038) := x"ffff";
    tmp(04039) := x"ffff";
    tmp(04040) := x"ffff";
    tmp(04041) := x"ffff";
    tmp(04042) := x"ffff";
    tmp(04043) := x"ffff";
    tmp(04044) := x"ffff";
    tmp(04045) := x"ffff";
    tmp(04046) := x"ffff";
    tmp(04047) := x"ffff";
    tmp(04048) := x"ffff";
    tmp(04049) := x"ffff";
    tmp(04050) := x"ffff";
    tmp(04051) := x"ffff";
    tmp(04052) := x"ffff";
    tmp(04053) := x"ffff";
    tmp(04054) := x"ffff";
    tmp(04055) := x"ffff";
    tmp(04056) := x"ffff";
    tmp(04057) := x"ffff";
    tmp(04058) := x"ffff";
    tmp(04059) := x"ffff";
    tmp(04060) := x"ffff";
    tmp(04061) := x"ffff";
    tmp(04062) := x"ffff";
    tmp(04063) := x"ffff";
    tmp(04064) := x"ffff";
    tmp(04065) := x"ffff";
    tmp(04066) := x"ffff";
    tmp(04067) := x"ffff";
    tmp(04068) := x"ffff";
    tmp(04069) := x"ffff";
    tmp(04070) := x"ffff";
    tmp(04071) := x"ffff";
    tmp(04072) := x"ffff";
    tmp(04073) := x"ffff";
    tmp(04074) := x"ffff";
    tmp(04075) := x"ffff";
    tmp(04076) := x"ffff";
    tmp(04077) := x"0820";
    tmp(04078) := x"0020";
    tmp(04079) := x"0020";
    tmp(04080) := x"0000";
    tmp(04081) := x"0020";
    tmp(04082) := x"0020";
    tmp(04083) := x"0020";
    tmp(04084) := x"0020";
    tmp(04085) := x"0020";
    tmp(04086) := x"0020";
    tmp(04087) := x"0020";
    tmp(04088) := x"0020";
    tmp(04089) := x"0020";
    tmp(04090) := x"0020";
    tmp(04091) := x"0040";
    tmp(04092) := x"0040";
    tmp(04093) := x"0040";
    tmp(04094) := x"0040";
    tmp(04095) := x"0040";
    tmp(04096) := x"0040";
    tmp(04097) := x"0040";
    tmp(04098) := x"0040";
    tmp(04099) := x"0040";
    tmp(04100) := x"0040";
    tmp(04101) := x"0040";
    tmp(04102) := x"0040";
    tmp(04103) := x"0840";
    tmp(04104) := x"0840";
    tmp(04105) := x"0040";
    tmp(04106) := x"0040";
    tmp(04107) := x"0040";
    tmp(04108) := x"0040";
    tmp(04109) := x"0040";
    tmp(04110) := x"0040";
    tmp(04111) := x"0040";
    tmp(04112) := x"0060";
    tmp(04113) := x"0040";
    tmp(04114) := x"0040";
    tmp(04115) := x"0040";
    tmp(04116) := x"0060";
    tmp(04117) := x"0060";
    tmp(04118) := x"0060";
    tmp(04119) := x"0060";
    tmp(04120) := x"0060";
    tmp(04121) := x"0060";
    tmp(04122) := x"0060";
    tmp(04123) := x"0060";
    tmp(04124) := x"0060";
    tmp(04125) := x"0060";
    tmp(04126) := x"0060";
    tmp(04127) := x"0060";
    tmp(04128) := x"0860";
    tmp(04129) := x"0860";
    tmp(04130) := x"0860";
    tmp(04131) := x"0860";
    tmp(04132) := x"0860";
    tmp(04133) := x"0860";
    tmp(04134) := x"0860";
    tmp(04135) := x"0860";
    tmp(04136) := x"0840";
    tmp(04137) := x"0840";
    tmp(04138) := x"0840";
    tmp(04139) := x"0840";
    tmp(04140) := x"0840";
    tmp(04141) := x"0840";
    tmp(04142) := x"0840";
    tmp(04143) := x"0840";
    tmp(04144) := x"0840";
    tmp(04145) := x"0820";
    tmp(04146) := x"0840";
    tmp(04147) := x"0840";
    tmp(04148) := x"0840";
    tmp(04149) := x"0820";
    tmp(04150) := x"0840";
    tmp(04151) := x"0840";
    tmp(04152) := x"0840";
    tmp(04153) := x"0840";
    tmp(04154) := x"0840";
    tmp(04155) := x"0840";
    tmp(04156) := x"0840";
    tmp(04157) := x"0840";
    tmp(04158) := x"0840";
    tmp(04159) := x"0840";
    tmp(04160) := x"0840";
    tmp(04161) := x"0840";
    tmp(04162) := x"0840";
    tmp(04163) := x"0840";
    tmp(04164) := x"0840";
    tmp(04165) := x"0840";
    tmp(04166) := x"0840";
    tmp(04167) := x"0840";
    tmp(04168) := x"0860";
    tmp(04169) := x"0860";
    tmp(04170) := x"0860";
    tmp(04171) := x"0860";
    tmp(04172) := x"0860";
    tmp(04173) := x"0860";
    tmp(04174) := x"0880";
    tmp(04175) := x"0880";
    tmp(04176) := x"0880";
    tmp(04177) := x"0880";
    tmp(04178) := x"0880";
    tmp(04179) := x"0880";
    tmp(04180) := x"0880";
    tmp(04181) := x"0880";
    tmp(04182) := x"0880";
    tmp(04183) := x"0880";
    tmp(04184) := x"08a0";
    tmp(04185) := x"0880";
    tmp(04186) := x"0860";
    tmp(04187) := x"0040";
    tmp(04188) := x"0020";
    tmp(04189) := x"0000";
    tmp(04190) := x"0000";
    tmp(04191) := x"0000";
    tmp(04192) := x"0000";
    tmp(04193) := x"0000";
    tmp(04194) := x"0000";
    tmp(04195) := x"0000";
    tmp(04196) := x"0000";
    tmp(04197) := x"0000";
    tmp(04198) := x"0000";
    tmp(04199) := x"0000";
    tmp(04200) := x"0000";
    tmp(04201) := x"0000";
    tmp(04202) := x"0000";
    tmp(04203) := x"0021";
    tmp(04204) := x"0841";
    tmp(04205) := x"0861";
    tmp(04206) := x"0882";
    tmp(04207) := x"10c3";
    tmp(04208) := x"1904";
    tmp(04209) := x"1943";
    tmp(04210) := x"1122";
    tmp(04211) := x"08c0";
    tmp(04212) := x"08a0";
    tmp(04213) := x"00a0";
    tmp(04214) := x"00a0";
    tmp(04215) := x"00a0";
    tmp(04216) := x"00a0";
    tmp(04217) := x"00a0";
    tmp(04218) := x"00a0";
    tmp(04219) := x"00a0";
    tmp(04220) := x"00c0";
    tmp(04221) := x"00c0";
    tmp(04222) := x"00a0";
    tmp(04223) := x"00c0";
    tmp(04224) := x"00a0";
    tmp(04225) := x"00c0";
    tmp(04226) := x"00c0";
    tmp(04227) := x"00c0";
    tmp(04228) := x"08c0";
    tmp(04229) := x"08c0";
    tmp(04230) := x"08c0";
    tmp(04231) := x"08c0";
    tmp(04232) := x"08c0";
    tmp(04233) := x"08c0";
    tmp(04234) := x"08c0";
    tmp(04235) := x"08c0";
    tmp(04236) := x"08c0";
    tmp(04237) := x"08c0";
    tmp(04238) := x"08c0";
    tmp(04239) := x"08c0";
    tmp(04240) := x"08c0";
    tmp(04241) := x"08c0";
    tmp(04242) := x"08c0";
    tmp(04243) := x"08c0";
    tmp(04244) := x"08c0";
    tmp(04245) := x"08c0";
    tmp(04246) := x"08c0";
    tmp(04247) := x"08c0";
    tmp(04248) := x"08c0";
    tmp(04249) := x"08c0";
    tmp(04250) := x"08c0";
    tmp(04251) := x"08c0";
    tmp(04252) := x"08c0";
    tmp(04253) := x"08c0";
    tmp(04254) := x"08c0";
    tmp(04255) := x"08c0";
    tmp(04256) := x"08c0";
    tmp(04257) := x"08c0";
    tmp(04258) := x"08c0";
    tmp(04259) := x"08c0";
    tmp(04260) := x"08c0";
    tmp(04261) := x"08c0";
    tmp(04262) := x"08c0";
    tmp(04263) := x"08c0";
    tmp(04264) := x"08c0";
    tmp(04265) := x"08c0";
    tmp(04266) := x"08c0";
    tmp(04267) := x"08c0";
    tmp(04268) := x"08c0";
    tmp(04269) := x"08a0";
    tmp(04270) := x"08a0";
    tmp(04271) := x"08a0";
    tmp(04272) := x"08a0";
    tmp(04273) := x"08a0";
    tmp(04274) := x"08a0";
    tmp(04275) := x"08a0";
    tmp(04276) := x"08a0";
    tmp(04277) := x"ffff";
    tmp(04278) := x"ffff";
    tmp(04279) := x"ffff";
    tmp(04280) := x"ffff";
    tmp(04281) := x"ffff";
    tmp(04282) := x"ffff";
    tmp(04283) := x"ffff";
    tmp(04284) := x"ffff";
    tmp(04285) := x"ffff";
    tmp(04286) := x"ffff";
    tmp(04287) := x"ffff";
    tmp(04288) := x"ffff";
    tmp(04289) := x"ffff";
    tmp(04290) := x"ffff";
    tmp(04291) := x"ffff";
    tmp(04292) := x"ffff";
    tmp(04293) := x"ffff";
    tmp(04294) := x"ffff";
    tmp(04295) := x"ffff";
    tmp(04296) := x"ffff";
    tmp(04297) := x"ffff";
    tmp(04298) := x"ffff";
    tmp(04299) := x"ffff";
    tmp(04300) := x"ffff";
    tmp(04301) := x"ffff";
    tmp(04302) := x"ffff";
    tmp(04303) := x"ffff";
    tmp(04304) := x"ffff";
    tmp(04305) := x"ffff";
    tmp(04306) := x"ffff";
    tmp(04307) := x"ffff";
    tmp(04308) := x"ffff";
    tmp(04309) := x"ffff";
    tmp(04310) := x"ffff";
    tmp(04311) := x"ffff";
    tmp(04312) := x"ffff";
    tmp(04313) := x"ffff";
    tmp(04314) := x"ffff";
    tmp(04315) := x"ffff";
    tmp(04316) := x"ffff";
    tmp(04317) := x"0020";
    tmp(04318) := x"0020";
    tmp(04319) := x"0020";
    tmp(04320) := x"0000";
    tmp(04321) := x"0020";
    tmp(04322) := x"0020";
    tmp(04323) := x"0020";
    tmp(04324) := x"0020";
    tmp(04325) := x"0020";
    tmp(04326) := x"0020";
    tmp(04327) := x"0020";
    tmp(04328) := x"0020";
    tmp(04329) := x"0020";
    tmp(04330) := x"0020";
    tmp(04331) := x"0040";
    tmp(04332) := x"0040";
    tmp(04333) := x"0040";
    tmp(04334) := x"0040";
    tmp(04335) := x"0040";
    tmp(04336) := x"0040";
    tmp(04337) := x"0040";
    tmp(04338) := x"0040";
    tmp(04339) := x"0040";
    tmp(04340) := x"0040";
    tmp(04341) := x"0040";
    tmp(04342) := x"0040";
    tmp(04343) := x"0040";
    tmp(04344) := x"0040";
    tmp(04345) := x"0040";
    tmp(04346) := x"0040";
    tmp(04347) := x"0040";
    tmp(04348) := x"0040";
    tmp(04349) := x"0040";
    tmp(04350) := x"0040";
    tmp(04351) := x"0040";
    tmp(04352) := x"0040";
    tmp(04353) := x"0040";
    tmp(04354) := x"0040";
    tmp(04355) := x"0040";
    tmp(04356) := x"0040";
    tmp(04357) := x"0040";
    tmp(04358) := x"0040";
    tmp(04359) := x"0060";
    tmp(04360) := x"0060";
    tmp(04361) := x"0060";
    tmp(04362) := x"0060";
    tmp(04363) := x"0060";
    tmp(04364) := x"0060";
    tmp(04365) := x"0060";
    tmp(04366) := x"0860";
    tmp(04367) := x"0860";
    tmp(04368) := x"0860";
    tmp(04369) := x"0860";
    tmp(04370) := x"0860";
    tmp(04371) := x"0860";
    tmp(04372) := x"0860";
    tmp(04373) := x"0860";
    tmp(04374) := x"0840";
    tmp(04375) := x"0840";
    tmp(04376) := x"0840";
    tmp(04377) := x"0840";
    tmp(04378) := x"0840";
    tmp(04379) := x"0840";
    tmp(04380) := x"0840";
    tmp(04381) := x"0840";
    tmp(04382) := x"0840";
    tmp(04383) := x"0840";
    tmp(04384) := x"0840";
    tmp(04385) := x"0840";
    tmp(04386) := x"0840";
    tmp(04387) := x"0840";
    tmp(04388) := x"0840";
    tmp(04389) := x"0840";
    tmp(04390) := x"0840";
    tmp(04391) := x"0840";
    tmp(04392) := x"0840";
    tmp(04393) := x"0840";
    tmp(04394) := x"0840";
    tmp(04395) := x"0840";
    tmp(04396) := x"0840";
    tmp(04397) := x"0840";
    tmp(04398) := x"0840";
    tmp(04399) := x"0840";
    tmp(04400) := x"0840";
    tmp(04401) := x"0840";
    tmp(04402) := x"0840";
    tmp(04403) := x"0840";
    tmp(04404) := x"0840";
    tmp(04405) := x"0840";
    tmp(04406) := x"0840";
    tmp(04407) := x"0840";
    tmp(04408) := x"0840";
    tmp(04409) := x"0860";
    tmp(04410) := x"0860";
    tmp(04411) := x"0860";
    tmp(04412) := x"0860";
    tmp(04413) := x"0860";
    tmp(04414) := x"0880";
    tmp(04415) := x"0880";
    tmp(04416) := x"0880";
    tmp(04417) := x"0880";
    tmp(04418) := x"0880";
    tmp(04419) := x"0880";
    tmp(04420) := x"0880";
    tmp(04421) := x"0880";
    tmp(04422) := x"0880";
    tmp(04423) := x"0880";
    tmp(04424) := x"0880";
    tmp(04425) := x"0880";
    tmp(04426) := x"08a0";
    tmp(04427) := x"08a0";
    tmp(04428) := x"08a0";
    tmp(04429) := x"0860";
    tmp(04430) := x"0040";
    tmp(04431) := x"0020";
    tmp(04432) := x"0000";
    tmp(04433) := x"0000";
    tmp(04434) := x"0000";
    tmp(04435) := x"0000";
    tmp(04436) := x"0000";
    tmp(04437) := x"0000";
    tmp(04438) := x"0000";
    tmp(04439) := x"0000";
    tmp(04440) := x"0000";
    tmp(04441) := x"0000";
    tmp(04442) := x"0000";
    tmp(04443) := x"0000";
    tmp(04444) := x"0000";
    tmp(04445) := x"0020";
    tmp(04446) := x"0841";
    tmp(04447) := x"0861";
    tmp(04448) := x"0882";
    tmp(04449) := x"10a3";
    tmp(04450) := x"1904";
    tmp(04451) := x"1923";
    tmp(04452) := x"1101";
    tmp(04453) := x"08a0";
    tmp(04454) := x"0080";
    tmp(04455) := x"00a0";
    tmp(04456) := x"00a0";
    tmp(04457) := x"00a0";
    tmp(04458) := x"00a0";
    tmp(04459) := x"00a0";
    tmp(04460) := x"00c0";
    tmp(04461) := x"00c0";
    tmp(04462) := x"00c0";
    tmp(04463) := x"00a0";
    tmp(04464) := x"00c0";
    tmp(04465) := x"00c0";
    tmp(04466) := x"00a0";
    tmp(04467) := x"08c0";
    tmp(04468) := x"08c0";
    tmp(04469) := x"08c0";
    tmp(04470) := x"08c0";
    tmp(04471) := x"08c0";
    tmp(04472) := x"08c0";
    tmp(04473) := x"08c0";
    tmp(04474) := x"08c0";
    tmp(04475) := x"08c0";
    tmp(04476) := x"08c0";
    tmp(04477) := x"08c0";
    tmp(04478) := x"08c0";
    tmp(04479) := x"08c0";
    tmp(04480) := x"08c0";
    tmp(04481) := x"08c0";
    tmp(04482) := x"08c0";
    tmp(04483) := x"08c0";
    tmp(04484) := x"08c0";
    tmp(04485) := x"08c0";
    tmp(04486) := x"08c0";
    tmp(04487) := x"08c0";
    tmp(04488) := x"08c0";
    tmp(04489) := x"08c0";
    tmp(04490) := x"08c0";
    tmp(04491) := x"08c0";
    tmp(04492) := x"08c0";
    tmp(04493) := x"08c0";
    tmp(04494) := x"08c0";
    tmp(04495) := x"08c0";
    tmp(04496) := x"08c0";
    tmp(04497) := x"08c0";
    tmp(04498) := x"08c0";
    tmp(04499) := x"08c0";
    tmp(04500) := x"08c0";
    tmp(04501) := x"08c0";
    tmp(04502) := x"08c0";
    tmp(04503) := x"08c0";
    tmp(04504) := x"08c0";
    tmp(04505) := x"08c0";
    tmp(04506) := x"08a0";
    tmp(04507) := x"08a0";
    tmp(04508) := x"08a0";
    tmp(04509) := x"08a0";
    tmp(04510) := x"08a0";
    tmp(04511) := x"08a0";
    tmp(04512) := x"08a0";
    tmp(04513) := x"08a0";
    tmp(04514) := x"08a0";
    tmp(04515) := x"08a0";
    tmp(04516) := x"08a0";
    tmp(04517) := x"ffff";
    tmp(04518) := x"ffff";
    tmp(04519) := x"ffff";
    tmp(04520) := x"ffff";
    tmp(04521) := x"ffff";
    tmp(04522) := x"ffff";
    tmp(04523) := x"ffff";
    tmp(04524) := x"ffff";
    tmp(04525) := x"ffff";
    tmp(04526) := x"ffff";
    tmp(04527) := x"ffff";
    tmp(04528) := x"ffff";
    tmp(04529) := x"ffff";
    tmp(04530) := x"ffff";
    tmp(04531) := x"ffff";
    tmp(04532) := x"ffff";
    tmp(04533) := x"ffff";
    tmp(04534) := x"ffff";
    tmp(04535) := x"ffff";
    tmp(04536) := x"ffff";
    tmp(04537) := x"ffff";
    tmp(04538) := x"ffff";
    tmp(04539) := x"ffff";
    tmp(04540) := x"ffff";
    tmp(04541) := x"ffff";
    tmp(04542) := x"ffff";
    tmp(04543) := x"ffff";
    tmp(04544) := x"ffff";
    tmp(04545) := x"ffff";
    tmp(04546) := x"ffff";
    tmp(04547) := x"ffff";
    tmp(04548) := x"ffff";
    tmp(04549) := x"ffff";
    tmp(04550) := x"ffff";
    tmp(04551) := x"ffff";
    tmp(04552) := x"ffff";
    tmp(04553) := x"ffff";
    tmp(04554) := x"ffff";
    tmp(04555) := x"ffff";
    tmp(04556) := x"ffff";
    tmp(04557) := x"0020";
    tmp(04558) := x"0020";
    tmp(04559) := x"0020";
    tmp(04560) := x"0000";
    tmp(04561) := x"0020";
    tmp(04562) := x"0020";
    tmp(04563) := x"0020";
    tmp(04564) := x"0020";
    tmp(04565) := x"0020";
    tmp(04566) := x"0020";
    tmp(04567) := x"0020";
    tmp(04568) := x"0020";
    tmp(04569) := x"0020";
    tmp(04570) := x"0020";
    tmp(04571) := x"0040";
    tmp(04572) := x"0040";
    tmp(04573) := x"0040";
    tmp(04574) := x"0040";
    tmp(04575) := x"0040";
    tmp(04576) := x"0040";
    tmp(04577) := x"0040";
    tmp(04578) := x"0040";
    tmp(04579) := x"0040";
    tmp(04580) := x"0040";
    tmp(04581) := x"0040";
    tmp(04582) := x"0040";
    tmp(04583) := x"0040";
    tmp(04584) := x"0040";
    tmp(04585) := x"0040";
    tmp(04586) := x"0040";
    tmp(04587) := x"0040";
    tmp(04588) := x"0040";
    tmp(04589) := x"0040";
    tmp(04590) := x"0040";
    tmp(04591) := x"0040";
    tmp(04592) := x"0040";
    tmp(04593) := x"0040";
    tmp(04594) := x"0040";
    tmp(04595) := x"0040";
    tmp(04596) := x"0040";
    tmp(04597) := x"0040";
    tmp(04598) := x"0040";
    tmp(04599) := x"0040";
    tmp(04600) := x"0040";
    tmp(04601) := x"0040";
    tmp(04602) := x"0060";
    tmp(04603) := x"0860";
    tmp(04604) := x"0860";
    tmp(04605) := x"0860";
    tmp(04606) := x"0860";
    tmp(04607) := x"0840";
    tmp(04608) := x"0860";
    tmp(04609) := x"0860";
    tmp(04610) := x"0840";
    tmp(04611) := x"0840";
    tmp(04612) := x"0840";
    tmp(04613) := x"0840";
    tmp(04614) := x"0840";
    tmp(04615) := x"0840";
    tmp(04616) := x"0840";
    tmp(04617) := x"0840";
    tmp(04618) := x"0840";
    tmp(04619) := x"0840";
    tmp(04620) := x"0840";
    tmp(04621) := x"0840";
    tmp(04622) := x"0840";
    tmp(04623) := x"0840";
    tmp(04624) := x"0840";
    tmp(04625) := x"0840";
    tmp(04626) := x"0840";
    tmp(04627) := x"0840";
    tmp(04628) := x"0820";
    tmp(04629) := x"0840";
    tmp(04630) := x"0840";
    tmp(04631) := x"0840";
    tmp(04632) := x"0840";
    tmp(04633) := x"0840";
    tmp(04634) := x"0840";
    tmp(04635) := x"0840";
    tmp(04636) := x"0840";
    tmp(04637) := x"0840";
    tmp(04638) := x"0840";
    tmp(04639) := x"0840";
    tmp(04640) := x"0840";
    tmp(04641) := x"0840";
    tmp(04642) := x"0840";
    tmp(04643) := x"0840";
    tmp(04644) := x"0840";
    tmp(04645) := x"0840";
    tmp(04646) := x"0840";
    tmp(04647) := x"0840";
    tmp(04648) := x"0860";
    tmp(04649) := x"0860";
    tmp(04650) := x"0860";
    tmp(04651) := x"0860";
    tmp(04652) := x"0860";
    tmp(04653) := x"0860";
    tmp(04654) := x"0860";
    tmp(04655) := x"0880";
    tmp(04656) := x"0880";
    tmp(04657) := x"0880";
    tmp(04658) := x"0880";
    tmp(04659) := x"0880";
    tmp(04660) := x"08a0";
    tmp(04661) := x"0880";
    tmp(04662) := x"0880";
    tmp(04663) := x"0880";
    tmp(04664) := x"0880";
    tmp(04665) := x"0880";
    tmp(04666) := x"0880";
    tmp(04667) := x"0880";
    tmp(04668) := x"08a0";
    tmp(04669) := x"08a0";
    tmp(04670) := x"08a0";
    tmp(04671) := x"0860";
    tmp(04672) := x"0040";
    tmp(04673) := x"0000";
    tmp(04674) := x"0000";
    tmp(04675) := x"0000";
    tmp(04676) := x"0000";
    tmp(04677) := x"0000";
    tmp(04678) := x"0000";
    tmp(04679) := x"0000";
    tmp(04680) := x"0000";
    tmp(04681) := x"0000";
    tmp(04682) := x"0000";
    tmp(04683) := x"0000";
    tmp(04684) := x"0000";
    tmp(04685) := x"0000";
    tmp(04686) := x"0000";
    tmp(04687) := x"0021";
    tmp(04688) := x"0841";
    tmp(04689) := x"0841";
    tmp(04690) := x"0862";
    tmp(04691) := x"1082";
    tmp(04692) := x"10a2";
    tmp(04693) := x"10c2";
    tmp(04694) := x"08c1";
    tmp(04695) := x"08a0";
    tmp(04696) := x"00a0";
    tmp(04697) := x"00a0";
    tmp(04698) := x"00a0";
    tmp(04699) := x"00a0";
    tmp(04700) := x"08a0";
    tmp(04701) := x"08a0";
    tmp(04702) := x"08a0";
    tmp(04703) := x"00a0";
    tmp(04704) := x"08a0";
    tmp(04705) := x"00c0";
    tmp(04706) := x"08c0";
    tmp(04707) := x"08c0";
    tmp(04708) := x"08c0";
    tmp(04709) := x"08c0";
    tmp(04710) := x"08c0";
    tmp(04711) := x"08c0";
    tmp(04712) := x"08c0";
    tmp(04713) := x"08c0";
    tmp(04714) := x"08c0";
    tmp(04715) := x"08c0";
    tmp(04716) := x"08c0";
    tmp(04717) := x"08c0";
    tmp(04718) := x"08c0";
    tmp(04719) := x"08c0";
    tmp(04720) := x"08c0";
    tmp(04721) := x"08c0";
    tmp(04722) := x"08c0";
    tmp(04723) := x"08c0";
    tmp(04724) := x"08c0";
    tmp(04725) := x"08c0";
    tmp(04726) := x"08c0";
    tmp(04727) := x"08c0";
    tmp(04728) := x"08c0";
    tmp(04729) := x"08c0";
    tmp(04730) := x"08c0";
    tmp(04731) := x"08c0";
    tmp(04732) := x"08c0";
    tmp(04733) := x"08c0";
    tmp(04734) := x"08c0";
    tmp(04735) := x"08c0";
    tmp(04736) := x"08c0";
    tmp(04737) := x"08c0";
    tmp(04738) := x"08c0";
    tmp(04739) := x"08c0";
    tmp(04740) := x"08c0";
    tmp(04741) := x"08c0";
    tmp(04742) := x"08c0";
    tmp(04743) := x"08c0";
    tmp(04744) := x"08c0";
    tmp(04745) := x"08c0";
    tmp(04746) := x"08c0";
    tmp(04747) := x"08a0";
    tmp(04748) := x"08a0";
    tmp(04749) := x"08a0";
    tmp(04750) := x"08a0";
    tmp(04751) := x"08a0";
    tmp(04752) := x"08a0";
    tmp(04753) := x"08a0";
    tmp(04754) := x"08a0";
    tmp(04755) := x"08a0";
    tmp(04756) := x"08a0";
    tmp(04757) := x"ffff";
    tmp(04758) := x"ffff";
    tmp(04759) := x"ffff";
    tmp(04760) := x"ffff";
    tmp(04761) := x"ffff";
    tmp(04762) := x"ffff";
    tmp(04763) := x"ffff";
    tmp(04764) := x"ffff";
    tmp(04765) := x"ffff";
    tmp(04766) := x"ffff";
    tmp(04767) := x"ffff";
    tmp(04768) := x"ffff";
    tmp(04769) := x"ffff";
    tmp(04770) := x"ffff";
    tmp(04771) := x"ffff";
    tmp(04772) := x"ffff";
    tmp(04773) := x"ffff";
    tmp(04774) := x"ffff";
    tmp(04775) := x"ffff";
    tmp(04776) := x"ffff";
    tmp(04777) := x"ffff";
    tmp(04778) := x"ffff";
    tmp(04779) := x"ffff";
    tmp(04780) := x"ffff";
    tmp(04781) := x"ffff";
    tmp(04782) := x"ffff";
    tmp(04783) := x"ffff";
    tmp(04784) := x"ffff";
    tmp(04785) := x"ffff";
    tmp(04786) := x"ffff";
    tmp(04787) := x"ffff";
    tmp(04788) := x"ffff";
    tmp(04789) := x"ffff";
    tmp(04790) := x"ffff";
    tmp(04791) := x"ffff";
    tmp(04792) := x"ffff";
    tmp(04793) := x"ffff";
    tmp(04794) := x"ffff";
    tmp(04795) := x"ffff";
    tmp(04796) := x"ffff";
    tmp(04797) := x"0020";
    tmp(04798) := x"0020";
    tmp(04799) := x"0820";
    tmp(04800) := x"0000";
    tmp(04801) := x"0020";
    tmp(04802) := x"0020";
    tmp(04803) := x"0020";
    tmp(04804) := x"0020";
    tmp(04805) := x"0020";
    tmp(04806) := x"0020";
    tmp(04807) := x"0020";
    tmp(04808) := x"0020";
    tmp(04809) := x"0020";
    tmp(04810) := x"0040";
    tmp(04811) := x"0040";
    tmp(04812) := x"0040";
    tmp(04813) := x"0040";
    tmp(04814) := x"0040";
    tmp(04815) := x"0040";
    tmp(04816) := x"0040";
    tmp(04817) := x"0040";
    tmp(04818) := x"0040";
    tmp(04819) := x"0040";
    tmp(04820) := x"0040";
    tmp(04821) := x"0040";
    tmp(04822) := x"0040";
    tmp(04823) := x"0040";
    tmp(04824) := x"0040";
    tmp(04825) := x"0040";
    tmp(04826) := x"0040";
    tmp(04827) := x"0040";
    tmp(04828) := x"0040";
    tmp(04829) := x"0040";
    tmp(04830) := x"0040";
    tmp(04831) := x"0040";
    tmp(04832) := x"0040";
    tmp(04833) := x"0040";
    tmp(04834) := x"0040";
    tmp(04835) := x"0040";
    tmp(04836) := x"0040";
    tmp(04837) := x"0040";
    tmp(04838) := x"0040";
    tmp(04839) := x"0040";
    tmp(04840) := x"0040";
    tmp(04841) := x"0840";
    tmp(04842) := x"0840";
    tmp(04843) := x"0840";
    tmp(04844) := x"0840";
    tmp(04845) := x"0840";
    tmp(04846) := x"0840";
    tmp(04847) := x"0840";
    tmp(04848) := x"0840";
    tmp(04849) := x"0840";
    tmp(04850) := x"0840";
    tmp(04851) := x"0840";
    tmp(04852) := x"0840";
    tmp(04853) := x"0840";
    tmp(04854) := x"0840";
    tmp(04855) := x"0840";
    tmp(04856) := x"0840";
    tmp(04857) := x"0840";
    tmp(04858) := x"0840";
    tmp(04859) := x"0840";
    tmp(04860) := x"0840";
    tmp(04861) := x"0840";
    tmp(04862) := x"0840";
    tmp(04863) := x"0840";
    tmp(04864) := x"0820";
    tmp(04865) := x"0840";
    tmp(04866) := x"0840";
    tmp(04867) := x"0840";
    tmp(04868) := x"0840";
    tmp(04869) := x"0840";
    tmp(04870) := x"0840";
    tmp(04871) := x"0840";
    tmp(04872) := x"0840";
    tmp(04873) := x"0840";
    tmp(04874) := x"0840";
    tmp(04875) := x"0840";
    tmp(04876) := x"0840";
    tmp(04877) := x"0840";
    tmp(04878) := x"0840";
    tmp(04879) := x"0840";
    tmp(04880) := x"0840";
    tmp(04881) := x"0840";
    tmp(04882) := x"0840";
    tmp(04883) := x"0840";
    tmp(04884) := x"0840";
    tmp(04885) := x"0840";
    tmp(04886) := x"0840";
    tmp(04887) := x"0840";
    tmp(04888) := x"0840";
    tmp(04889) := x"0860";
    tmp(04890) := x"0860";
    tmp(04891) := x"0860";
    tmp(04892) := x"0860";
    tmp(04893) := x"0860";
    tmp(04894) := x"0880";
    tmp(04895) := x"0880";
    tmp(04896) := x"0880";
    tmp(04897) := x"0880";
    tmp(04898) := x"0880";
    tmp(04899) := x"0880";
    tmp(04900) := x"0880";
    tmp(04901) := x"0880";
    tmp(04902) := x"0880";
    tmp(04903) := x"0880";
    tmp(04904) := x"0880";
    tmp(04905) := x"0880";
    tmp(04906) := x"0880";
    tmp(04907) := x"0880";
    tmp(04908) := x"0880";
    tmp(04909) := x"0880";
    tmp(04910) := x"0880";
    tmp(04911) := x"0880";
    tmp(04912) := x"0880";
    tmp(04913) := x"0860";
    tmp(04914) := x"0020";
    tmp(04915) := x"0000";
    tmp(04916) := x"0000";
    tmp(04917) := x"0000";
    tmp(04918) := x"0000";
    tmp(04919) := x"0000";
    tmp(04920) := x"0000";
    tmp(04921) := x"0000";
    tmp(04922) := x"0000";
    tmp(04923) := x"0000";
    tmp(04924) := x"0000";
    tmp(04925) := x"0000";
    tmp(04926) := x"0000";
    tmp(04927) := x"0000";
    tmp(04928) := x"0020";
    tmp(04929) := x"0021";
    tmp(04930) := x"0841";
    tmp(04931) := x"0841";
    tmp(04932) := x"0841";
    tmp(04933) := x"0841";
    tmp(04934) := x"0881";
    tmp(04935) := x"08a1";
    tmp(04936) := x"08a0";
    tmp(04937) := x"00a0";
    tmp(04938) := x"00a0";
    tmp(04939) := x"00a0";
    tmp(04940) := x"08a0";
    tmp(04941) := x"08a0";
    tmp(04942) := x"08a0";
    tmp(04943) := x"08a0";
    tmp(04944) := x"08a0";
    tmp(04945) := x"08c0";
    tmp(04946) := x"08c0";
    tmp(04947) := x"08c0";
    tmp(04948) := x"08c0";
    tmp(04949) := x"08c0";
    tmp(04950) := x"08c0";
    tmp(04951) := x"08c0";
    tmp(04952) := x"08c0";
    tmp(04953) := x"08c0";
    tmp(04954) := x"08c0";
    tmp(04955) := x"08c0";
    tmp(04956) := x"08c0";
    tmp(04957) := x"08c0";
    tmp(04958) := x"08c0";
    tmp(04959) := x"08c0";
    tmp(04960) := x"08c0";
    tmp(04961) := x"08c0";
    tmp(04962) := x"08c0";
    tmp(04963) := x"08c0";
    tmp(04964) := x"08c0";
    tmp(04965) := x"08c0";
    tmp(04966) := x"08c0";
    tmp(04967) := x"08c0";
    tmp(04968) := x"08c0";
    tmp(04969) := x"08c0";
    tmp(04970) := x"08c0";
    tmp(04971) := x"08c0";
    tmp(04972) := x"08c0";
    tmp(04973) := x"08c0";
    tmp(04974) := x"08c0";
    tmp(04975) := x"08c0";
    tmp(04976) := x"08c0";
    tmp(04977) := x"08c0";
    tmp(04978) := x"08c0";
    tmp(04979) := x"08c0";
    tmp(04980) := x"08c0";
    tmp(04981) := x"08c0";
    tmp(04982) := x"08c0";
    tmp(04983) := x"08c0";
    tmp(04984) := x"08c0";
    tmp(04985) := x"08c0";
    tmp(04986) := x"08c0";
    tmp(04987) := x"08a0";
    tmp(04988) := x"08a0";
    tmp(04989) := x"08a0";
    tmp(04990) := x"08a0";
    tmp(04991) := x"08a0";
    tmp(04992) := x"08a0";
    tmp(04993) := x"08a0";
    tmp(04994) := x"08a0";
    tmp(04995) := x"08a0";
    tmp(04996) := x"08a0";
    tmp(04997) := x"ffff";
    tmp(04998) := x"ffff";
    tmp(04999) := x"ffff";
    tmp(05000) := x"ffff";
    tmp(05001) := x"ffff";
    tmp(05002) := x"ffff";
    tmp(05003) := x"ffff";
    tmp(05004) := x"ffff";
    tmp(05005) := x"ffff";
    tmp(05006) := x"ffff";
    tmp(05007) := x"ffff";
    tmp(05008) := x"ffff";
    tmp(05009) := x"ffff";
    tmp(05010) := x"ffff";
    tmp(05011) := x"ffff";
    tmp(05012) := x"ffff";
    tmp(05013) := x"ffff";
    tmp(05014) := x"ffff";
    tmp(05015) := x"ffff";
    tmp(05016) := x"ffff";
    tmp(05017) := x"ffff";
    tmp(05018) := x"ffff";
    tmp(05019) := x"ffff";
    tmp(05020) := x"ffff";
    tmp(05021) := x"ffff";
    tmp(05022) := x"ffff";
    tmp(05023) := x"ffff";
    tmp(05024) := x"ffff";
    tmp(05025) := x"ffff";
    tmp(05026) := x"ffff";
    tmp(05027) := x"ffff";
    tmp(05028) := x"ffff";
    tmp(05029) := x"ffff";
    tmp(05030) := x"ffff";
    tmp(05031) := x"ffff";
    tmp(05032) := x"ffff";
    tmp(05033) := x"ffff";
    tmp(05034) := x"ffff";
    tmp(05035) := x"ffff";
    tmp(05036) := x"ffff";
    tmp(05037) := x"0820";
    tmp(05038) := x"0020";
    tmp(05039) := x"0020";
    tmp(05040) := x"0000";
    tmp(05041) := x"0020";
    tmp(05042) := x"0020";
    tmp(05043) := x"0020";
    tmp(05044) := x"0020";
    tmp(05045) := x"0020";
    tmp(05046) := x"0020";
    tmp(05047) := x"0020";
    tmp(05048) := x"0020";
    tmp(05049) := x"0020";
    tmp(05050) := x"0040";
    tmp(05051) := x"0040";
    tmp(05052) := x"0040";
    tmp(05053) := x"0040";
    tmp(05054) := x"0040";
    tmp(05055) := x"0040";
    tmp(05056) := x"0040";
    tmp(05057) := x"0040";
    tmp(05058) := x"0040";
    tmp(05059) := x"0040";
    tmp(05060) := x"0040";
    tmp(05061) := x"0040";
    tmp(05062) := x"0040";
    tmp(05063) := x"0040";
    tmp(05064) := x"0040";
    tmp(05065) := x"0040";
    tmp(05066) := x"0040";
    tmp(05067) := x"0040";
    tmp(05068) := x"0040";
    tmp(05069) := x"0040";
    tmp(05070) := x"0040";
    tmp(05071) := x"0040";
    tmp(05072) := x"0040";
    tmp(05073) := x"0040";
    tmp(05074) := x"0040";
    tmp(05075) := x"0040";
    tmp(05076) := x"0040";
    tmp(05077) := x"0040";
    tmp(05078) := x"0040";
    tmp(05079) := x"0040";
    tmp(05080) := x"0840";
    tmp(05081) := x"0840";
    tmp(05082) := x"0840";
    tmp(05083) := x"0840";
    tmp(05084) := x"0840";
    tmp(05085) := x"0840";
    tmp(05086) := x"0840";
    tmp(05087) := x"0840";
    tmp(05088) := x"0840";
    tmp(05089) := x"0840";
    tmp(05090) := x"0840";
    tmp(05091) := x"0840";
    tmp(05092) := x"0840";
    tmp(05093) := x"0840";
    tmp(05094) := x"0840";
    tmp(05095) := x"0840";
    tmp(05096) := x"0840";
    tmp(05097) := x"0840";
    tmp(05098) := x"0840";
    tmp(05099) := x"0840";
    tmp(05100) := x"0840";
    tmp(05101) := x"0840";
    tmp(05102) := x"0840";
    tmp(05103) := x"0840";
    tmp(05104) := x"0840";
    tmp(05105) := x"0840";
    tmp(05106) := x"0840";
    tmp(05107) := x"0840";
    tmp(05108) := x"0840";
    tmp(05109) := x"0840";
    tmp(05110) := x"0840";
    tmp(05111) := x"0840";
    tmp(05112) := x"0840";
    tmp(05113) := x"0840";
    tmp(05114) := x"0840";
    tmp(05115) := x"0840";
    tmp(05116) := x"0840";
    tmp(05117) := x"0840";
    tmp(05118) := x"0840";
    tmp(05119) := x"0840";
    tmp(05120) := x"0840";
    tmp(05121) := x"0840";
    tmp(05122) := x"0840";
    tmp(05123) := x"0840";
    tmp(05124) := x"0840";
    tmp(05125) := x"0840";
    tmp(05126) := x"0840";
    tmp(05127) := x"0860";
    tmp(05128) := x"0860";
    tmp(05129) := x"0860";
    tmp(05130) := x"0860";
    tmp(05131) := x"0860";
    tmp(05132) := x"0860";
    tmp(05133) := x"0860";
    tmp(05134) := x"0880";
    tmp(05135) := x"0880";
    tmp(05136) := x"0880";
    tmp(05137) := x"0880";
    tmp(05138) := x"0880";
    tmp(05139) := x"0880";
    tmp(05140) := x"0880";
    tmp(05141) := x"0880";
    tmp(05142) := x"08a0";
    tmp(05143) := x"0880";
    tmp(05144) := x"0880";
    tmp(05145) := x"0880";
    tmp(05146) := x"0880";
    tmp(05147) := x"0880";
    tmp(05148) := x"08a0";
    tmp(05149) := x"0880";
    tmp(05150) := x"0880";
    tmp(05151) := x"0880";
    tmp(05152) := x"0880";
    tmp(05153) := x"0880";
    tmp(05154) := x"0860";
    tmp(05155) := x"0840";
    tmp(05156) := x"0000";
    tmp(05157) := x"0000";
    tmp(05158) := x"0000";
    tmp(05159) := x"0000";
    tmp(05160) := x"0000";
    tmp(05161) := x"0000";
    tmp(05162) := x"0000";
    tmp(05163) := x"0000";
    tmp(05164) := x"0000";
    tmp(05165) := x"0000";
    tmp(05166) := x"0000";
    tmp(05167) := x"0000";
    tmp(05168) := x"0000";
    tmp(05169) := x"0000";
    tmp(05170) := x"0021";
    tmp(05171) := x"0841";
    tmp(05172) := x"0841";
    tmp(05173) := x"0821";
    tmp(05174) := x"0841";
    tmp(05175) := x"0841";
    tmp(05176) := x"0881";
    tmp(05177) := x"08a0";
    tmp(05178) := x"0880";
    tmp(05179) := x"08a0";
    tmp(05180) := x"08a0";
    tmp(05181) := x"08a0";
    tmp(05182) := x"08a0";
    tmp(05183) := x"08a0";
    tmp(05184) := x"08a0";
    tmp(05185) := x"08a0";
    tmp(05186) := x"08a0";
    tmp(05187) := x"08a0";
    tmp(05188) := x"08c0";
    tmp(05189) := x"08c0";
    tmp(05190) := x"08c0";
    tmp(05191) := x"08c0";
    tmp(05192) := x"08c0";
    tmp(05193) := x"08c0";
    tmp(05194) := x"08c0";
    tmp(05195) := x"08c0";
    tmp(05196) := x"08c0";
    tmp(05197) := x"08c0";
    tmp(05198) := x"08c0";
    tmp(05199) := x"08c0";
    tmp(05200) := x"08c0";
    tmp(05201) := x"08c0";
    tmp(05202) := x"08e0";
    tmp(05203) := x"08e0";
    tmp(05204) := x"08c0";
    tmp(05205) := x"08c0";
    tmp(05206) := x"08c0";
    tmp(05207) := x"08e0";
    tmp(05208) := x"08e0";
    tmp(05209) := x"08c0";
    tmp(05210) := x"08e0";
    tmp(05211) := x"08c0";
    tmp(05212) := x"08c0";
    tmp(05213) := x"08c0";
    tmp(05214) := x"08c0";
    tmp(05215) := x"08c0";
    tmp(05216) := x"08c0";
    tmp(05217) := x"08c0";
    tmp(05218) := x"08c0";
    tmp(05219) := x"08c0";
    tmp(05220) := x"08c0";
    tmp(05221) := x"08c0";
    tmp(05222) := x"08c0";
    tmp(05223) := x"08c0";
    tmp(05224) := x"08c0";
    tmp(05225) := x"08c0";
    tmp(05226) := x"08c0";
    tmp(05227) := x"08c0";
    tmp(05228) := x"08c0";
    tmp(05229) := x"08a0";
    tmp(05230) := x"08a0";
    tmp(05231) := x"08a0";
    tmp(05232) := x"08a0";
    tmp(05233) := x"08a0";
    tmp(05234) := x"08a0";
    tmp(05235) := x"08a0";
    tmp(05236) := x"08a0";
    tmp(05237) := x"ffff";
    tmp(05238) := x"ffff";
    tmp(05239) := x"ffff";
    tmp(05240) := x"ffff";
    tmp(05241) := x"ffff";
    tmp(05242) := x"ffff";
    tmp(05243) := x"ffff";
    tmp(05244) := x"ffff";
    tmp(05245) := x"ffff";
    tmp(05246) := x"ffff";
    tmp(05247) := x"ffff";
    tmp(05248) := x"ffff";
    tmp(05249) := x"ffff";
    tmp(05250) := x"ffff";
    tmp(05251) := x"ffff";
    tmp(05252) := x"ffff";
    tmp(05253) := x"ffff";
    tmp(05254) := x"ffff";
    tmp(05255) := x"ffff";
    tmp(05256) := x"ffff";
    tmp(05257) := x"ffff";
    tmp(05258) := x"ffff";
    tmp(05259) := x"ffff";
    tmp(05260) := x"ffff";
    tmp(05261) := x"ffff";
    tmp(05262) := x"ffff";
    tmp(05263) := x"ffff";
    tmp(05264) := x"ffff";
    tmp(05265) := x"ffff";
    tmp(05266) := x"ffff";
    tmp(05267) := x"ffff";
    tmp(05268) := x"ffff";
    tmp(05269) := x"ffff";
    tmp(05270) := x"ffff";
    tmp(05271) := x"ffff";
    tmp(05272) := x"ffff";
    tmp(05273) := x"ffff";
    tmp(05274) := x"ffff";
    tmp(05275) := x"ffff";
    tmp(05276) := x"ffff";
    tmp(05277) := x"0820";
    tmp(05278) := x"0820";
    tmp(05279) := x"0020";
    tmp(05280) := x"0000";
    tmp(05281) := x"0020";
    tmp(05282) := x"0020";
    tmp(05283) := x"0020";
    tmp(05284) := x"0020";
    tmp(05285) := x"0020";
    tmp(05286) := x"0020";
    tmp(05287) := x"0020";
    tmp(05288) := x"0020";
    tmp(05289) := x"0020";
    tmp(05290) := x"0040";
    tmp(05291) := x"0040";
    tmp(05292) := x"0040";
    tmp(05293) := x"0040";
    tmp(05294) := x"0040";
    tmp(05295) := x"0040";
    tmp(05296) := x"0040";
    tmp(05297) := x"0040";
    tmp(05298) := x"0040";
    tmp(05299) := x"0040";
    tmp(05300) := x"0040";
    tmp(05301) := x"0040";
    tmp(05302) := x"0040";
    tmp(05303) := x"0040";
    tmp(05304) := x"0040";
    tmp(05305) := x"0040";
    tmp(05306) := x"0040";
    tmp(05307) := x"0040";
    tmp(05308) := x"0040";
    tmp(05309) := x"0020";
    tmp(05310) := x"0020";
    tmp(05311) := x"0020";
    tmp(05312) := x"0020";
    tmp(05313) := x"0040";
    tmp(05314) := x"0040";
    tmp(05315) := x"0040";
    tmp(05316) := x"0040";
    tmp(05317) := x"0040";
    tmp(05318) := x"0840";
    tmp(05319) := x"0840";
    tmp(05320) := x"0840";
    tmp(05321) := x"0840";
    tmp(05322) := x"0840";
    tmp(05323) := x"0840";
    tmp(05324) := x"0840";
    tmp(05325) := x"0840";
    tmp(05326) := x"0840";
    tmp(05327) := x"0840";
    tmp(05328) := x"0840";
    tmp(05329) := x"0840";
    tmp(05330) := x"0840";
    tmp(05331) := x"0840";
    tmp(05332) := x"0840";
    tmp(05333) := x"0840";
    tmp(05334) := x"0840";
    tmp(05335) := x"0840";
    tmp(05336) := x"0840";
    tmp(05337) := x"0840";
    tmp(05338) := x"0840";
    tmp(05339) := x"0840";
    tmp(05340) := x"0840";
    tmp(05341) := x"0840";
    tmp(05342) := x"0840";
    tmp(05343) := x"0840";
    tmp(05344) := x"0840";
    tmp(05345) := x"0840";
    tmp(05346) := x"0840";
    tmp(05347) := x"0840";
    tmp(05348) := x"0840";
    tmp(05349) := x"0840";
    tmp(05350) := x"0840";
    tmp(05351) := x"0840";
    tmp(05352) := x"0840";
    tmp(05353) := x"0840";
    tmp(05354) := x"0840";
    tmp(05355) := x"0840";
    tmp(05356) := x"0840";
    tmp(05357) := x"0840";
    tmp(05358) := x"0840";
    tmp(05359) := x"0840";
    tmp(05360) := x"0840";
    tmp(05361) := x"0840";
    tmp(05362) := x"0840";
    tmp(05363) := x"0840";
    tmp(05364) := x"0840";
    tmp(05365) := x"0840";
    tmp(05366) := x"0840";
    tmp(05367) := x"0860";
    tmp(05368) := x"0860";
    tmp(05369) := x"0860";
    tmp(05370) := x"0860";
    tmp(05371) := x"0860";
    tmp(05372) := x"0860";
    tmp(05373) := x"0860";
    tmp(05374) := x"0880";
    tmp(05375) := x"0880";
    tmp(05376) := x"0880";
    tmp(05377) := x"0880";
    tmp(05378) := x"0880";
    tmp(05379) := x"0880";
    tmp(05380) := x"0880";
    tmp(05381) := x"0880";
    tmp(05382) := x"0880";
    tmp(05383) := x"0880";
    tmp(05384) := x"0880";
    tmp(05385) := x"0880";
    tmp(05386) := x"0880";
    tmp(05387) := x"0880";
    tmp(05388) := x"0880";
    tmp(05389) := x"0880";
    tmp(05390) := x"0880";
    tmp(05391) := x"0880";
    tmp(05392) := x"0860";
    tmp(05393) := x"0840";
    tmp(05394) := x"0860";
    tmp(05395) := x"0880";
    tmp(05396) := x"0880";
    tmp(05397) := x"0020";
    tmp(05398) := x"0000";
    tmp(05399) := x"0000";
    tmp(05400) := x"0000";
    tmp(05401) := x"0000";
    tmp(05402) := x"0000";
    tmp(05403) := x"0000";
    tmp(05404) := x"0000";
    tmp(05405) := x"0000";
    tmp(05406) := x"0000";
    tmp(05407) := x"0000";
    tmp(05408) := x"0000";
    tmp(05409) := x"0000";
    tmp(05410) := x"0000";
    tmp(05411) := x"0020";
    tmp(05412) := x"0021";
    tmp(05413) := x"0821";
    tmp(05414) := x"0021";
    tmp(05415) := x"0021";
    tmp(05416) := x"0021";
    tmp(05417) := x"0861";
    tmp(05418) := x"08a1";
    tmp(05419) := x"0880";
    tmp(05420) := x"08a0";
    tmp(05421) := x"00a0";
    tmp(05422) := x"08a0";
    tmp(05423) := x"08a0";
    tmp(05424) := x"08a0";
    tmp(05425) := x"08a0";
    tmp(05426) := x"08a0";
    tmp(05427) := x"08a0";
    tmp(05428) := x"08c0";
    tmp(05429) := x"00a0";
    tmp(05430) := x"08c0";
    tmp(05431) := x"08c0";
    tmp(05432) := x"08a0";
    tmp(05433) := x"08c0";
    tmp(05434) := x"08a0";
    tmp(05435) := x"08c0";
    tmp(05436) := x"08c0";
    tmp(05437) := x"08c0";
    tmp(05438) := x"08c0";
    tmp(05439) := x"08c0";
    tmp(05440) := x"08c0";
    tmp(05441) := x"08c0";
    tmp(05442) := x"08c0";
    tmp(05443) := x"08e0";
    tmp(05444) := x"08e0";
    tmp(05445) := x"08c0";
    tmp(05446) := x"08e0";
    tmp(05447) := x"08c0";
    tmp(05448) := x"08e0";
    tmp(05449) := x"08c0";
    tmp(05450) := x"08c0";
    tmp(05451) := x"08e0";
    tmp(05452) := x"08e0";
    tmp(05453) := x"08e0";
    tmp(05454) := x"08e0";
    tmp(05455) := x"08c0";
    tmp(05456) := x"08c0";
    tmp(05457) := x"08e0";
    tmp(05458) := x"08e0";
    tmp(05459) := x"08c0";
    tmp(05460) := x"08e0";
    tmp(05461) := x"08c0";
    tmp(05462) := x"08c0";
    tmp(05463) := x"08c0";
    tmp(05464) := x"08e0";
    tmp(05465) := x"08c0";
    tmp(05466) := x"08c0";
    tmp(05467) := x"08c0";
    tmp(05468) := x"08c0";
    tmp(05469) := x"08c0";
    tmp(05470) := x"08a0";
    tmp(05471) := x"08a0";
    tmp(05472) := x"08a0";
    tmp(05473) := x"08a0";
    tmp(05474) := x"08a0";
    tmp(05475) := x"08a0";
    tmp(05476) := x"08a0";
    tmp(05477) := x"ffff";
    tmp(05478) := x"ffff";
    tmp(05479) := x"ffff";
    tmp(05480) := x"ffff";
    tmp(05481) := x"ffff";
    tmp(05482) := x"ffff";
    tmp(05483) := x"ffff";
    tmp(05484) := x"ffff";
    tmp(05485) := x"ffff";
    tmp(05486) := x"ffff";
    tmp(05487) := x"ffff";
    tmp(05488) := x"ffff";
    tmp(05489) := x"ffff";
    tmp(05490) := x"ffff";
    tmp(05491) := x"ffff";
    tmp(05492) := x"ffff";
    tmp(05493) := x"ffff";
    tmp(05494) := x"ffff";
    tmp(05495) := x"ffff";
    tmp(05496) := x"ffff";
    tmp(05497) := x"ffff";
    tmp(05498) := x"ffff";
    tmp(05499) := x"ffff";
    tmp(05500) := x"ffff";
    tmp(05501) := x"ffff";
    tmp(05502) := x"ffff";
    tmp(05503) := x"ffff";
    tmp(05504) := x"ffff";
    tmp(05505) := x"ffff";
    tmp(05506) := x"ffff";
    tmp(05507) := x"ffff";
    tmp(05508) := x"ffff";
    tmp(05509) := x"ffff";
    tmp(05510) := x"ffff";
    tmp(05511) := x"ffff";
    tmp(05512) := x"ffff";
    tmp(05513) := x"ffff";
    tmp(05514) := x"ffff";
    tmp(05515) := x"ffff";
    tmp(05516) := x"ffff";
    tmp(05517) := x"0820";
    tmp(05518) := x"0820";
    tmp(05519) := x"0820";
    tmp(05520) := x"0000";
    tmp(05521) := x"0020";
    tmp(05522) := x"0020";
    tmp(05523) := x"0020";
    tmp(05524) := x"0020";
    tmp(05525) := x"0020";
    tmp(05526) := x"0020";
    tmp(05527) := x"0020";
    tmp(05528) := x"0020";
    tmp(05529) := x"0040";
    tmp(05530) := x"0040";
    tmp(05531) := x"0040";
    tmp(05532) := x"0040";
    tmp(05533) := x"0040";
    tmp(05534) := x"0040";
    tmp(05535) := x"0040";
    tmp(05536) := x"0040";
    tmp(05537) := x"0040";
    tmp(05538) := x"0040";
    tmp(05539) := x"0040";
    tmp(05540) := x"0040";
    tmp(05541) := x"0040";
    tmp(05542) := x"0040";
    tmp(05543) := x"0040";
    tmp(05544) := x"0040";
    tmp(05545) := x"0040";
    tmp(05546) := x"0040";
    tmp(05547) := x"0020";
    tmp(05548) := x"0020";
    tmp(05549) := x"0020";
    tmp(05550) := x"0020";
    tmp(05551) := x"0020";
    tmp(05552) := x"0020";
    tmp(05553) := x"0020";
    tmp(05554) := x"0020";
    tmp(05555) := x"0020";
    tmp(05556) := x"0040";
    tmp(05557) := x"0840";
    tmp(05558) := x"0840";
    tmp(05559) := x"0840";
    tmp(05560) := x"0840";
    tmp(05561) := x"0840";
    tmp(05562) := x"0840";
    tmp(05563) := x"0840";
    tmp(05564) := x"0840";
    tmp(05565) := x"0840";
    tmp(05566) := x"0840";
    tmp(05567) := x"0840";
    tmp(05568) := x"0840";
    tmp(05569) := x"0840";
    tmp(05570) := x"0840";
    tmp(05571) := x"0840";
    tmp(05572) := x"0840";
    tmp(05573) := x"0840";
    tmp(05574) := x"0840";
    tmp(05575) := x"0840";
    tmp(05576) := x"0840";
    tmp(05577) := x"0840";
    tmp(05578) := x"0840";
    tmp(05579) := x"0840";
    tmp(05580) := x"0840";
    tmp(05581) := x"0840";
    tmp(05582) := x"0840";
    tmp(05583) := x"0840";
    tmp(05584) := x"0840";
    tmp(05585) := x"0840";
    tmp(05586) := x"0840";
    tmp(05587) := x"0840";
    tmp(05588) := x"0840";
    tmp(05589) := x"0840";
    tmp(05590) := x"0840";
    tmp(05591) := x"0840";
    tmp(05592) := x"0840";
    tmp(05593) := x"0840";
    tmp(05594) := x"0840";
    tmp(05595) := x"0840";
    tmp(05596) := x"0840";
    tmp(05597) := x"0840";
    tmp(05598) := x"0840";
    tmp(05599) := x"0840";
    tmp(05600) := x"0840";
    tmp(05601) := x"0840";
    tmp(05602) := x"0840";
    tmp(05603) := x"0840";
    tmp(05604) := x"0840";
    tmp(05605) := x"0840";
    tmp(05606) := x"0860";
    tmp(05607) := x"0860";
    tmp(05608) := x"0860";
    tmp(05609) := x"0860";
    tmp(05610) := x"0860";
    tmp(05611) := x"0860";
    tmp(05612) := x"0860";
    tmp(05613) := x"0860";
    tmp(05614) := x"0860";
    tmp(05615) := x"0880";
    tmp(05616) := x"0880";
    tmp(05617) := x"0880";
    tmp(05618) := x"0880";
    tmp(05619) := x"0880";
    tmp(05620) := x"0880";
    tmp(05621) := x"0880";
    tmp(05622) := x"0880";
    tmp(05623) := x"0880";
    tmp(05624) := x"0880";
    tmp(05625) := x"0880";
    tmp(05626) := x"0880";
    tmp(05627) := x"08a0";
    tmp(05628) := x"0880";
    tmp(05629) := x"08a0";
    tmp(05630) := x"08a0";
    tmp(05631) := x"0840";
    tmp(05632) := x"0020";
    tmp(05633) := x"0840";
    tmp(05634) := x"0860";
    tmp(05635) := x"0880";
    tmp(05636) := x"0880";
    tmp(05637) := x"0880";
    tmp(05638) := x"0040";
    tmp(05639) := x"0000";
    tmp(05640) := x"0000";
    tmp(05641) := x"0000";
    tmp(05642) := x"0000";
    tmp(05643) := x"0000";
    tmp(05644) := x"0000";
    tmp(05645) := x"0000";
    tmp(05646) := x"0000";
    tmp(05647) := x"0000";
    tmp(05648) := x"0000";
    tmp(05649) := x"0000";
    tmp(05650) := x"0000";
    tmp(05651) := x"0000";
    tmp(05652) := x"0020";
    tmp(05653) := x"0021";
    tmp(05654) := x"0841";
    tmp(05655) := x"0021";
    tmp(05656) := x"0021";
    tmp(05657) := x"0021";
    tmp(05658) := x"0841";
    tmp(05659) := x"08a1";
    tmp(05660) := x"0880";
    tmp(05661) := x"08a0";
    tmp(05662) := x"08a0";
    tmp(05663) := x"08a0";
    tmp(05664) := x"08a0";
    tmp(05665) := x"08a0";
    tmp(05666) := x"08a0";
    tmp(05667) := x"08a0";
    tmp(05668) := x"08a0";
    tmp(05669) := x"08a0";
    tmp(05670) := x"08a0";
    tmp(05671) := x"08a0";
    tmp(05672) := x"08a0";
    tmp(05673) := x"08a0";
    tmp(05674) := x"08a0";
    tmp(05675) := x"08a0";
    tmp(05676) := x"08c0";
    tmp(05677) := x"08c0";
    tmp(05678) := x"08c0";
    tmp(05679) := x"08c0";
    tmp(05680) := x"08c0";
    tmp(05681) := x"08c0";
    tmp(05682) := x"08c0";
    tmp(05683) := x"08c0";
    tmp(05684) := x"08c0";
    tmp(05685) := x"08c0";
    tmp(05686) := x"08c0";
    tmp(05687) := x"08c0";
    tmp(05688) := x"08e0";
    tmp(05689) := x"08c0";
    tmp(05690) := x"08e0";
    tmp(05691) := x"08c0";
    tmp(05692) := x"08e0";
    tmp(05693) := x"08e0";
    tmp(05694) := x"08e0";
    tmp(05695) := x"08e0";
    tmp(05696) := x"08e0";
    tmp(05697) := x"08e0";
    tmp(05698) := x"08c0";
    tmp(05699) := x"08c0";
    tmp(05700) := x"08e0";
    tmp(05701) := x"08e0";
    tmp(05702) := x"08c0";
    tmp(05703) := x"08c0";
    tmp(05704) := x"08e0";
    tmp(05705) := x"08c0";
    tmp(05706) := x"08c0";
    tmp(05707) := x"08c0";
    tmp(05708) := x"08c0";
    tmp(05709) := x"08c0";
    tmp(05710) := x"08c0";
    tmp(05711) := x"08c0";
    tmp(05712) := x"08c0";
    tmp(05713) := x"08a0";
    tmp(05714) := x"08a0";
    tmp(05715) := x"08a0";
    tmp(05716) := x"08a0";
    tmp(05717) := x"ffff";
    tmp(05718) := x"ffff";
    tmp(05719) := x"ffff";
    tmp(05720) := x"ffff";
    tmp(05721) := x"ffff";
    tmp(05722) := x"ffff";
    tmp(05723) := x"ffff";
    tmp(05724) := x"ffff";
    tmp(05725) := x"ffff";
    tmp(05726) := x"ffff";
    tmp(05727) := x"ffff";
    tmp(05728) := x"ffff";
    tmp(05729) := x"ffff";
    tmp(05730) := x"ffff";
    tmp(05731) := x"ffff";
    tmp(05732) := x"ffff";
    tmp(05733) := x"ffff";
    tmp(05734) := x"ffff";
    tmp(05735) := x"ffff";
    tmp(05736) := x"ffff";
    tmp(05737) := x"ffff";
    tmp(05738) := x"ffff";
    tmp(05739) := x"ffff";
    tmp(05740) := x"ffff";
    tmp(05741) := x"ffff";
    tmp(05742) := x"ffff";
    tmp(05743) := x"ffff";
    tmp(05744) := x"ffff";
    tmp(05745) := x"ffff";
    tmp(05746) := x"ffff";
    tmp(05747) := x"ffff";
    tmp(05748) := x"ffff";
    tmp(05749) := x"ffff";
    tmp(05750) := x"ffff";
    tmp(05751) := x"ffff";
    tmp(05752) := x"ffff";
    tmp(05753) := x"ffff";
    tmp(05754) := x"ffff";
    tmp(05755) := x"ffff";
    tmp(05756) := x"ffff";
    tmp(05757) := x"0820";
    tmp(05758) := x"0820";
    tmp(05759) := x"0820";
    tmp(05760) := x"0000";
    tmp(05761) := x"0020";
    tmp(05762) := x"0020";
    tmp(05763) := x"0020";
    tmp(05764) := x"0020";
    tmp(05765) := x"0020";
    tmp(05766) := x"0020";
    tmp(05767) := x"0040";
    tmp(05768) := x"0040";
    tmp(05769) := x"0040";
    tmp(05770) := x"0040";
    tmp(05771) := x"0040";
    tmp(05772) := x"0040";
    tmp(05773) := x"0040";
    tmp(05774) := x"0040";
    tmp(05775) := x"0040";
    tmp(05776) := x"0040";
    tmp(05777) := x"0040";
    tmp(05778) := x"0040";
    tmp(05779) := x"0040";
    tmp(05780) := x"0040";
    tmp(05781) := x"0040";
    tmp(05782) := x"0040";
    tmp(05783) := x"0040";
    tmp(05784) := x"0020";
    tmp(05785) := x"0020";
    tmp(05786) := x"0020";
    tmp(05787) := x"0020";
    tmp(05788) := x"0020";
    tmp(05789) := x"0020";
    tmp(05790) := x"0020";
    tmp(05791) := x"0020";
    tmp(05792) := x"0020";
    tmp(05793) := x"0020";
    tmp(05794) := x"0020";
    tmp(05795) := x"0820";
    tmp(05796) := x"0820";
    tmp(05797) := x"0820";
    tmp(05798) := x"0820";
    tmp(05799) := x"0820";
    tmp(05800) := x"0820";
    tmp(05801) := x"0840";
    tmp(05802) := x"0840";
    tmp(05803) := x"0840";
    tmp(05804) := x"0840";
    tmp(05805) := x"0840";
    tmp(05806) := x"0840";
    tmp(05807) := x"0840";
    tmp(05808) := x"0840";
    tmp(05809) := x"0840";
    tmp(05810) := x"0840";
    tmp(05811) := x"0840";
    tmp(05812) := x"0840";
    tmp(05813) := x"0840";
    tmp(05814) := x"0840";
    tmp(05815) := x"0840";
    tmp(05816) := x"0840";
    tmp(05817) := x"0840";
    tmp(05818) := x"0840";
    tmp(05819) := x"0840";
    tmp(05820) := x"0840";
    tmp(05821) := x"0840";
    tmp(05822) := x"0840";
    tmp(05823) := x"0840";
    tmp(05824) := x"0840";
    tmp(05825) := x"0840";
    tmp(05826) := x"0840";
    tmp(05827) := x"0840";
    tmp(05828) := x"0840";
    tmp(05829) := x"0840";
    tmp(05830) := x"0840";
    tmp(05831) := x"0840";
    tmp(05832) := x"0840";
    tmp(05833) := x"0840";
    tmp(05834) := x"0840";
    tmp(05835) := x"0840";
    tmp(05836) := x"0840";
    tmp(05837) := x"0840";
    tmp(05838) := x"0840";
    tmp(05839) := x"0840";
    tmp(05840) := x"0840";
    tmp(05841) := x"0840";
    tmp(05842) := x"0840";
    tmp(05843) := x"0840";
    tmp(05844) := x"0840";
    tmp(05845) := x"0840";
    tmp(05846) := x"0860";
    tmp(05847) := x"0860";
    tmp(05848) := x"0860";
    tmp(05849) := x"0860";
    tmp(05850) := x"0860";
    tmp(05851) := x"0860";
    tmp(05852) := x"0860";
    tmp(05853) := x"0860";
    tmp(05854) := x"0860";
    tmp(05855) := x"0880";
    tmp(05856) := x"0880";
    tmp(05857) := x"0880";
    tmp(05858) := x"0880";
    tmp(05859) := x"0880";
    tmp(05860) := x"08a0";
    tmp(05861) := x"0880";
    tmp(05862) := x"0880";
    tmp(05863) := x"0880";
    tmp(05864) := x"0880";
    tmp(05865) := x"0880";
    tmp(05866) := x"0880";
    tmp(05867) := x"0880";
    tmp(05868) := x"0880";
    tmp(05869) := x"0880";
    tmp(05870) := x"0040";
    tmp(05871) := x"0000";
    tmp(05872) := x"0000";
    tmp(05873) := x"0840";
    tmp(05874) := x"0860";
    tmp(05875) := x"0880";
    tmp(05876) := x"0880";
    tmp(05877) := x"0880";
    tmp(05878) := x"0880";
    tmp(05879) := x"0860";
    tmp(05880) := x"0000";
    tmp(05881) := x"0000";
    tmp(05882) := x"0000";
    tmp(05883) := x"0000";
    tmp(05884) := x"0000";
    tmp(05885) := x"0000";
    tmp(05886) := x"0000";
    tmp(05887) := x"0000";
    tmp(05888) := x"0000";
    tmp(05889) := x"0000";
    tmp(05890) := x"0000";
    tmp(05891) := x"0000";
    tmp(05892) := x"0000";
    tmp(05893) := x"0020";
    tmp(05894) := x"0821";
    tmp(05895) := x"0841";
    tmp(05896) := x"0021";
    tmp(05897) := x"0021";
    tmp(05898) := x"0020";
    tmp(05899) := x"0841";
    tmp(05900) := x"08a1";
    tmp(05901) := x"0880";
    tmp(05902) := x"0880";
    tmp(05903) := x"0880";
    tmp(05904) := x"0880";
    tmp(05905) := x"08a0";
    tmp(05906) := x"08a0";
    tmp(05907) := x"08a0";
    tmp(05908) := x"08a0";
    tmp(05909) := x"08a0";
    tmp(05910) := x"08a0";
    tmp(05911) := x"08a0";
    tmp(05912) := x"08a0";
    tmp(05913) := x"08a0";
    tmp(05914) := x"08a0";
    tmp(05915) := x"08a0";
    tmp(05916) := x"08a0";
    tmp(05917) := x"08a0";
    tmp(05918) := x"08a0";
    tmp(05919) := x"08c0";
    tmp(05920) := x"08c0";
    tmp(05921) := x"08c0";
    tmp(05922) := x"08c0";
    tmp(05923) := x"08c0";
    tmp(05924) := x"08c0";
    tmp(05925) := x"08c0";
    tmp(05926) := x"08c0";
    tmp(05927) := x"08c0";
    tmp(05928) := x"08c0";
    tmp(05929) := x"08c0";
    tmp(05930) := x"08c0";
    tmp(05931) := x"08e0";
    tmp(05932) := x"08c0";
    tmp(05933) := x"08c0";
    tmp(05934) := x"08e0";
    tmp(05935) := x"08c0";
    tmp(05936) := x"08e0";
    tmp(05937) := x"08c0";
    tmp(05938) := x"08c0";
    tmp(05939) := x"08c0";
    tmp(05940) := x"08c0";
    tmp(05941) := x"08e0";
    tmp(05942) := x"08c0";
    tmp(05943) := x"08e0";
    tmp(05944) := x"08c0";
    tmp(05945) := x"08e0";
    tmp(05946) := x"08c0";
    tmp(05947) := x"08c0";
    tmp(05948) := x"08c0";
    tmp(05949) := x"08c0";
    tmp(05950) := x"08c0";
    tmp(05951) := x"08c0";
    tmp(05952) := x"08a0";
    tmp(05953) := x"08a0";
    tmp(05954) := x"08a0";
    tmp(05955) := x"08a0";
    tmp(05956) := x"08a0";
    tmp(05957) := x"ffff";
    tmp(05958) := x"ffff";
    tmp(05959) := x"ffff";
    tmp(05960) := x"ffff";
    tmp(05961) := x"ffff";
    tmp(05962) := x"ffff";
    tmp(05963) := x"ffff";
    tmp(05964) := x"ffff";
    tmp(05965) := x"ffff";
    tmp(05966) := x"ffff";
    tmp(05967) := x"ffff";
    tmp(05968) := x"ffff";
    tmp(05969) := x"ffff";
    tmp(05970) := x"ffff";
    tmp(05971) := x"ffff";
    tmp(05972) := x"ffff";
    tmp(05973) := x"ffff";
    tmp(05974) := x"ffff";
    tmp(05975) := x"ffff";
    tmp(05976) := x"ffff";
    tmp(05977) := x"ffff";
    tmp(05978) := x"ffff";
    tmp(05979) := x"ffff";
    tmp(05980) := x"ffff";
    tmp(05981) := x"ffff";
    tmp(05982) := x"ffff";
    tmp(05983) := x"ffff";
    tmp(05984) := x"ffff";
    tmp(05985) := x"ffff";
    tmp(05986) := x"ffff";
    tmp(05987) := x"ffff";
    tmp(05988) := x"ffff";
    tmp(05989) := x"ffff";
    tmp(05990) := x"ffff";
    tmp(05991) := x"ffff";
    tmp(05992) := x"ffff";
    tmp(05993) := x"ffff";
    tmp(05994) := x"ffff";
    tmp(05995) := x"ffff";
    tmp(05996) := x"ffff";
    tmp(05997) := x"0820";
    tmp(05998) := x"0820";
    tmp(05999) := x"0020";
    tmp(06000) := x"0000";
    tmp(06001) := x"0020";
    tmp(06002) := x"0020";
    tmp(06003) := x"0020";
    tmp(06004) := x"0020";
    tmp(06005) := x"0020";
    tmp(06006) := x"0020";
    tmp(06007) := x"0040";
    tmp(06008) := x"0040";
    tmp(06009) := x"0040";
    tmp(06010) := x"0040";
    tmp(06011) := x"0040";
    tmp(06012) := x"0040";
    tmp(06013) := x"0040";
    tmp(06014) := x"0040";
    tmp(06015) := x"0040";
    tmp(06016) := x"0040";
    tmp(06017) := x"0840";
    tmp(06018) := x"0040";
    tmp(06019) := x"0040";
    tmp(06020) := x"0840";
    tmp(06021) := x"0840";
    tmp(06022) := x"0040";
    tmp(06023) := x"0020";
    tmp(06024) := x"0020";
    tmp(06025) := x"0020";
    tmp(06026) := x"0020";
    tmp(06027) := x"0020";
    tmp(06028) := x"0020";
    tmp(06029) := x"0020";
    tmp(06030) := x"0020";
    tmp(06031) := x"0020";
    tmp(06032) := x"0020";
    tmp(06033) := x"0020";
    tmp(06034) := x"0820";
    tmp(06035) := x"0820";
    tmp(06036) := x"0820";
    tmp(06037) := x"0820";
    tmp(06038) := x"0820";
    tmp(06039) := x"0820";
    tmp(06040) := x"0820";
    tmp(06041) := x"0820";
    tmp(06042) := x"0820";
    tmp(06043) := x"0840";
    tmp(06044) := x"0840";
    tmp(06045) := x"0840";
    tmp(06046) := x"0840";
    tmp(06047) := x"0840";
    tmp(06048) := x"0840";
    tmp(06049) := x"0840";
    tmp(06050) := x"0840";
    tmp(06051) := x"0840";
    tmp(06052) := x"0840";
    tmp(06053) := x"0840";
    tmp(06054) := x"0840";
    tmp(06055) := x"0840";
    tmp(06056) := x"0840";
    tmp(06057) := x"0840";
    tmp(06058) := x"0840";
    tmp(06059) := x"0840";
    tmp(06060) := x"0840";
    tmp(06061) := x"0840";
    tmp(06062) := x"0840";
    tmp(06063) := x"0840";
    tmp(06064) := x"0840";
    tmp(06065) := x"0840";
    tmp(06066) := x"0840";
    tmp(06067) := x"0840";
    tmp(06068) := x"0840";
    tmp(06069) := x"0840";
    tmp(06070) := x"0840";
    tmp(06071) := x"0840";
    tmp(06072) := x"0840";
    tmp(06073) := x"0840";
    tmp(06074) := x"0840";
    tmp(06075) := x"0840";
    tmp(06076) := x"0840";
    tmp(06077) := x"0840";
    tmp(06078) := x"0840";
    tmp(06079) := x"0840";
    tmp(06080) := x"0840";
    tmp(06081) := x"0840";
    tmp(06082) := x"0840";
    tmp(06083) := x"0840";
    tmp(06084) := x"0840";
    tmp(06085) := x"0840";
    tmp(06086) := x"0860";
    tmp(06087) := x"0860";
    tmp(06088) := x"0860";
    tmp(06089) := x"0860";
    tmp(06090) := x"0860";
    tmp(06091) := x"0860";
    tmp(06092) := x"0860";
    tmp(06093) := x"0860";
    tmp(06094) := x"0880";
    tmp(06095) := x"0880";
    tmp(06096) := x"0880";
    tmp(06097) := x"0880";
    tmp(06098) := x"0880";
    tmp(06099) := x"0880";
    tmp(06100) := x"0880";
    tmp(06101) := x"08a0";
    tmp(06102) := x"0880";
    tmp(06103) := x"0880";
    tmp(06104) := x"08a0";
    tmp(06105) := x"0880";
    tmp(06106) := x"0880";
    tmp(06107) := x"08a0";
    tmp(06108) := x"0880";
    tmp(06109) := x"0020";
    tmp(06110) := x"0000";
    tmp(06111) := x"0000";
    tmp(06112) := x"0000";
    tmp(06113) := x"0840";
    tmp(06114) := x"0880";
    tmp(06115) := x"0880";
    tmp(06116) := x"0880";
    tmp(06117) := x"0880";
    tmp(06118) := x"0880";
    tmp(06119) := x"0880";
    tmp(06120) := x"0860";
    tmp(06121) := x"0000";
    tmp(06122) := x"0000";
    tmp(06123) := x"0000";
    tmp(06124) := x"0000";
    tmp(06125) := x"0000";
    tmp(06126) := x"0000";
    tmp(06127) := x"0000";
    tmp(06128) := x"0000";
    tmp(06129) := x"0000";
    tmp(06130) := x"0000";
    tmp(06131) := x"0000";
    tmp(06132) := x"0000";
    tmp(06133) := x"0000";
    tmp(06134) := x"0020";
    tmp(06135) := x"0821";
    tmp(06136) := x"0841";
    tmp(06137) := x"0841";
    tmp(06138) := x"0021";
    tmp(06139) := x"0020";
    tmp(06140) := x"0841";
    tmp(06141) := x"0881";
    tmp(06142) := x"0880";
    tmp(06143) := x"0880";
    tmp(06144) := x"0880";
    tmp(06145) := x"0880";
    tmp(06146) := x"0880";
    tmp(06147) := x"0880";
    tmp(06148) := x"0880";
    tmp(06149) := x"0880";
    tmp(06150) := x"0880";
    tmp(06151) := x"0880";
    tmp(06152) := x"0880";
    tmp(06153) := x"0880";
    tmp(06154) := x"0880";
    tmp(06155) := x"08a0";
    tmp(06156) := x"08a0";
    tmp(06157) := x"08a0";
    tmp(06158) := x"08a0";
    tmp(06159) := x"08a0";
    tmp(06160) := x"08a0";
    tmp(06161) := x"08a0";
    tmp(06162) := x"08a0";
    tmp(06163) := x"08c0";
    tmp(06164) := x"08c0";
    tmp(06165) := x"08a0";
    tmp(06166) := x"08c0";
    tmp(06167) := x"08c0";
    tmp(06168) := x"08c0";
    tmp(06169) := x"08c0";
    tmp(06170) := x"08c0";
    tmp(06171) := x"08c0";
    tmp(06172) := x"08c0";
    tmp(06173) := x"08c0";
    tmp(06174) := x"08c0";
    tmp(06175) := x"08c0";
    tmp(06176) := x"08c0";
    tmp(06177) := x"08c0";
    tmp(06178) := x"08c0";
    tmp(06179) := x"08c0";
    tmp(06180) := x"08c0";
    tmp(06181) := x"08c0";
    tmp(06182) := x"08e0";
    tmp(06183) := x"08c0";
    tmp(06184) := x"08c0";
    tmp(06185) := x"08c0";
    tmp(06186) := x"08c0";
    tmp(06187) := x"08c0";
    tmp(06188) := x"08c0";
    tmp(06189) := x"08c0";
    tmp(06190) := x"08c0";
    tmp(06191) := x"08a0";
    tmp(06192) := x"08a0";
    tmp(06193) := x"08a0";
    tmp(06194) := x"08a0";
    tmp(06195) := x"08a0";
    tmp(06196) := x"08a0";
    tmp(06197) := x"ffff";
    tmp(06198) := x"ffff";
    tmp(06199) := x"ffff";
    tmp(06200) := x"ffff";
    tmp(06201) := x"ffff";
    tmp(06202) := x"ffff";
    tmp(06203) := x"ffff";
    tmp(06204) := x"ffff";
    tmp(06205) := x"ffff";
    tmp(06206) := x"ffff";
    tmp(06207) := x"ffff";
    tmp(06208) := x"ffff";
    tmp(06209) := x"ffff";
    tmp(06210) := x"ffff";
    tmp(06211) := x"ffff";
    tmp(06212) := x"ffff";
    tmp(06213) := x"ffff";
    tmp(06214) := x"ffff";
    tmp(06215) := x"ffff";
    tmp(06216) := x"ffff";
    tmp(06217) := x"ffff";
    tmp(06218) := x"ffff";
    tmp(06219) := x"ffff";
    tmp(06220) := x"ffff";
    tmp(06221) := x"ffff";
    tmp(06222) := x"ffff";
    tmp(06223) := x"ffff";
    tmp(06224) := x"ffff";
    tmp(06225) := x"ffff";
    tmp(06226) := x"ffff";
    tmp(06227) := x"ffff";
    tmp(06228) := x"ffff";
    tmp(06229) := x"ffff";
    tmp(06230) := x"ffff";
    tmp(06231) := x"ffff";
    tmp(06232) := x"ffff";
    tmp(06233) := x"ffff";
    tmp(06234) := x"ffff";
    tmp(06235) := x"ffff";
    tmp(06236) := x"ffff";
    tmp(06237) := x"0820";
    tmp(06238) := x"0820";
    tmp(06239) := x"0820";
    tmp(06240) := x"0000";
    tmp(06241) := x"0020";
    tmp(06242) := x"0020";
    tmp(06243) := x"0020";
    tmp(06244) := x"0020";
    tmp(06245) := x"0020";
    tmp(06246) := x"0040";
    tmp(06247) := x"0040";
    tmp(06248) := x"0040";
    tmp(06249) := x"0040";
    tmp(06250) := x"0040";
    tmp(06251) := x"0040";
    tmp(06252) := x"0040";
    tmp(06253) := x"0040";
    tmp(06254) := x"0040";
    tmp(06255) := x"0040";
    tmp(06256) := x"0040";
    tmp(06257) := x"0840";
    tmp(06258) := x"0040";
    tmp(06259) := x"0840";
    tmp(06260) := x"0840";
    tmp(06261) := x"0820";
    tmp(06262) := x"0820";
    tmp(06263) := x"0820";
    tmp(06264) := x"0020";
    tmp(06265) := x"0020";
    tmp(06266) := x"0020";
    tmp(06267) := x"0020";
    tmp(06268) := x"0020";
    tmp(06269) := x"0020";
    tmp(06270) := x"0020";
    tmp(06271) := x"0020";
    tmp(06272) := x"0820";
    tmp(06273) := x"0820";
    tmp(06274) := x"0820";
    tmp(06275) := x"0820";
    tmp(06276) := x"0820";
    tmp(06277) := x"0820";
    tmp(06278) := x"0820";
    tmp(06279) := x"0820";
    tmp(06280) := x"0820";
    tmp(06281) := x"0820";
    tmp(06282) := x"0820";
    tmp(06283) := x"0820";
    tmp(06284) := x"0820";
    tmp(06285) := x"0820";
    tmp(06286) := x"0840";
    tmp(06287) := x"0840";
    tmp(06288) := x"0840";
    tmp(06289) := x"0840";
    tmp(06290) := x"0840";
    tmp(06291) := x"0840";
    tmp(06292) := x"0840";
    tmp(06293) := x"0840";
    tmp(06294) := x"0840";
    tmp(06295) := x"0840";
    tmp(06296) := x"0840";
    tmp(06297) := x"0840";
    tmp(06298) := x"0840";
    tmp(06299) := x"0840";
    tmp(06300) := x"0840";
    tmp(06301) := x"0840";
    tmp(06302) := x"0840";
    tmp(06303) := x"0840";
    tmp(06304) := x"0840";
    tmp(06305) := x"0840";
    tmp(06306) := x"0840";
    tmp(06307) := x"0840";
    tmp(06308) := x"0840";
    tmp(06309) := x"0840";
    tmp(06310) := x"0840";
    tmp(06311) := x"0840";
    tmp(06312) := x"0840";
    tmp(06313) := x"0840";
    tmp(06314) := x"0840";
    tmp(06315) := x"0840";
    tmp(06316) := x"0840";
    tmp(06317) := x"0840";
    tmp(06318) := x"0840";
    tmp(06319) := x"0840";
    tmp(06320) := x"0840";
    tmp(06321) := x"0840";
    tmp(06322) := x"0840";
    tmp(06323) := x"0840";
    tmp(06324) := x"0840";
    tmp(06325) := x"0860";
    tmp(06326) := x"0860";
    tmp(06327) := x"0860";
    tmp(06328) := x"0860";
    tmp(06329) := x"0860";
    tmp(06330) := x"0860";
    tmp(06331) := x"0860";
    tmp(06332) := x"0860";
    tmp(06333) := x"0860";
    tmp(06334) := x"0880";
    tmp(06335) := x"0880";
    tmp(06336) := x"0880";
    tmp(06337) := x"0880";
    tmp(06338) := x"0880";
    tmp(06339) := x"0880";
    tmp(06340) := x"08a0";
    tmp(06341) := x"08a0";
    tmp(06342) := x"08a0";
    tmp(06343) := x"08a0";
    tmp(06344) := x"08a0";
    tmp(06345) := x"08a0";
    tmp(06346) := x"08a0";
    tmp(06347) := x"0860";
    tmp(06348) := x"0020";
    tmp(06349) := x"0000";
    tmp(06350) := x"0000";
    tmp(06351) := x"0000";
    tmp(06352) := x"0000";
    tmp(06353) := x"0841";
    tmp(06354) := x"0881";
    tmp(06355) := x"0880";
    tmp(06356) := x"0880";
    tmp(06357) := x"0880";
    tmp(06358) := x"0880";
    tmp(06359) := x"0880";
    tmp(06360) := x"0880";
    tmp(06361) := x"0860";
    tmp(06362) := x"0000";
    tmp(06363) := x"0000";
    tmp(06364) := x"0000";
    tmp(06365) := x"0000";
    tmp(06366) := x"0000";
    tmp(06367) := x"0000";
    tmp(06368) := x"0000";
    tmp(06369) := x"0000";
    tmp(06370) := x"0000";
    tmp(06371) := x"0000";
    tmp(06372) := x"0000";
    tmp(06373) := x"0000";
    tmp(06374) := x"0000";
    tmp(06375) := x"0020";
    tmp(06376) := x"0821";
    tmp(06377) := x"0841";
    tmp(06378) := x"0821";
    tmp(06379) := x"0021";
    tmp(06380) := x"0020";
    tmp(06381) := x"0841";
    tmp(06382) := x"0881";
    tmp(06383) := x"0880";
    tmp(06384) := x"0880";
    tmp(06385) := x"0880";
    tmp(06386) := x"0880";
    tmp(06387) := x"0880";
    tmp(06388) := x"0880";
    tmp(06389) := x"0880";
    tmp(06390) := x"0880";
    tmp(06391) := x"0880";
    tmp(06392) := x"0880";
    tmp(06393) := x"0880";
    tmp(06394) := x"0880";
    tmp(06395) := x"0880";
    tmp(06396) := x"0880";
    tmp(06397) := x"0880";
    tmp(06398) := x"0880";
    tmp(06399) := x"08a0";
    tmp(06400) := x"0880";
    tmp(06401) := x"08a0";
    tmp(06402) := x"08a0";
    tmp(06403) := x"08a0";
    tmp(06404) := x"08a0";
    tmp(06405) := x"08a0";
    tmp(06406) := x"08a0";
    tmp(06407) := x"08a0";
    tmp(06408) := x"08a0";
    tmp(06409) := x"08a0";
    tmp(06410) := x"08a0";
    tmp(06411) := x"08c0";
    tmp(06412) := x"08c0";
    tmp(06413) := x"08c0";
    tmp(06414) := x"08c0";
    tmp(06415) := x"08c0";
    tmp(06416) := x"08c0";
    tmp(06417) := x"08c0";
    tmp(06418) := x"08c0";
    tmp(06419) := x"08c0";
    tmp(06420) := x"08c0";
    tmp(06421) := x"08c0";
    tmp(06422) := x"08c0";
    tmp(06423) := x"08c0";
    tmp(06424) := x"08c0";
    tmp(06425) := x"08c0";
    tmp(06426) := x"08c0";
    tmp(06427) := x"08c0";
    tmp(06428) := x"08c0";
    tmp(06429) := x"08c0";
    tmp(06430) := x"08c0";
    tmp(06431) := x"08c0";
    tmp(06432) := x"08c0";
    tmp(06433) := x"08a0";
    tmp(06434) := x"08a0";
    tmp(06435) := x"08a0";
    tmp(06436) := x"08a0";
    tmp(06437) := x"ffff";
    tmp(06438) := x"ffff";
    tmp(06439) := x"ffff";
    tmp(06440) := x"ffff";
    tmp(06441) := x"ffff";
    tmp(06442) := x"ffff";
    tmp(06443) := x"ffff";
    tmp(06444) := x"ffff";
    tmp(06445) := x"ffff";
    tmp(06446) := x"ffff";
    tmp(06447) := x"ffff";
    tmp(06448) := x"ffff";
    tmp(06449) := x"ffff";
    tmp(06450) := x"ffff";
    tmp(06451) := x"ffff";
    tmp(06452) := x"ffff";
    tmp(06453) := x"ffff";
    tmp(06454) := x"ffff";
    tmp(06455) := x"ffff";
    tmp(06456) := x"ffff";
    tmp(06457) := x"ffff";
    tmp(06458) := x"ffff";
    tmp(06459) := x"ffff";
    tmp(06460) := x"ffff";
    tmp(06461) := x"ffff";
    tmp(06462) := x"ffff";
    tmp(06463) := x"ffff";
    tmp(06464) := x"ffff";
    tmp(06465) := x"ffff";
    tmp(06466) := x"ffff";
    tmp(06467) := x"ffff";
    tmp(06468) := x"ffff";
    tmp(06469) := x"ffff";
    tmp(06470) := x"ffff";
    tmp(06471) := x"ffff";
    tmp(06472) := x"ffff";
    tmp(06473) := x"ffff";
    tmp(06474) := x"ffff";
    tmp(06475) := x"ffff";
    tmp(06476) := x"ffff";
    tmp(06477) := x"0820";
    tmp(06478) := x"0820";
    tmp(06479) := x"0820";
    tmp(06480) := x"0000";
    tmp(06481) := x"0020";
    tmp(06482) := x"0020";
    tmp(06483) := x"0020";
    tmp(06484) := x"0020";
    tmp(06485) := x"0040";
    tmp(06486) := x"0040";
    tmp(06487) := x"0040";
    tmp(06488) := x"0040";
    tmp(06489) := x"0040";
    tmp(06490) := x"0040";
    tmp(06491) := x"0040";
    tmp(06492) := x"0040";
    tmp(06493) := x"0040";
    tmp(06494) := x"0840";
    tmp(06495) := x"0840";
    tmp(06496) := x"0840";
    tmp(06497) := x"0840";
    tmp(06498) := x"0840";
    tmp(06499) := x"0840";
    tmp(06500) := x"0820";
    tmp(06501) := x"0820";
    tmp(06502) := x"0820";
    tmp(06503) := x"0820";
    tmp(06504) := x"0820";
    tmp(06505) := x"0820";
    tmp(06506) := x"0820";
    tmp(06507) := x"0020";
    tmp(06508) := x"0820";
    tmp(06509) := x"0820";
    tmp(06510) := x"0820";
    tmp(06511) := x"0820";
    tmp(06512) := x"0820";
    tmp(06513) := x"0820";
    tmp(06514) := x"0820";
    tmp(06515) := x"0820";
    tmp(06516) := x"0820";
    tmp(06517) := x"0820";
    tmp(06518) := x"0820";
    tmp(06519) := x"0820";
    tmp(06520) := x"0820";
    tmp(06521) := x"0820";
    tmp(06522) := x"0820";
    tmp(06523) := x"0820";
    tmp(06524) := x"0840";
    tmp(06525) := x"0840";
    tmp(06526) := x"0840";
    tmp(06527) := x"0840";
    tmp(06528) := x"0840";
    tmp(06529) := x"0840";
    tmp(06530) := x"0840";
    tmp(06531) := x"0840";
    tmp(06532) := x"0840";
    tmp(06533) := x"0840";
    tmp(06534) := x"0840";
    tmp(06535) := x"0840";
    tmp(06536) := x"0840";
    tmp(06537) := x"0840";
    tmp(06538) := x"0840";
    tmp(06539) := x"0841";
    tmp(06540) := x"0840";
    tmp(06541) := x"0840";
    tmp(06542) := x"0840";
    tmp(06543) := x"0840";
    tmp(06544) := x"0840";
    tmp(06545) := x"0840";
    tmp(06546) := x"0840";
    tmp(06547) := x"0840";
    tmp(06548) := x"0840";
    tmp(06549) := x"0840";
    tmp(06550) := x"0840";
    tmp(06551) := x"0840";
    tmp(06552) := x"0840";
    tmp(06553) := x"0840";
    tmp(06554) := x"0840";
    tmp(06555) := x"0840";
    tmp(06556) := x"0840";
    tmp(06557) := x"0840";
    tmp(06558) := x"0840";
    tmp(06559) := x"0840";
    tmp(06560) := x"0840";
    tmp(06561) := x"0840";
    tmp(06562) := x"0840";
    tmp(06563) := x"0840";
    tmp(06564) := x"0840";
    tmp(06565) := x"0860";
    tmp(06566) := x"0860";
    tmp(06567) := x"0860";
    tmp(06568) := x"0860";
    tmp(06569) := x"0860";
    tmp(06570) := x"0860";
    tmp(06571) := x"0860";
    tmp(06572) := x"0860";
    tmp(06573) := x"0860";
    tmp(06574) := x"0880";
    tmp(06575) := x"0880";
    tmp(06576) := x"0880";
    tmp(06577) := x"0880";
    tmp(06578) := x"0880";
    tmp(06579) := x"0880";
    tmp(06580) := x"08a0";
    tmp(06581) := x"08a0";
    tmp(06582) := x"08a0";
    tmp(06583) := x"0880";
    tmp(06584) := x"0880";
    tmp(06585) := x"0880";
    tmp(06586) := x"0860";
    tmp(06587) := x"0020";
    tmp(06588) := x"0000";
    tmp(06589) := x"0000";
    tmp(06590) := x"0000";
    tmp(06591) := x"0000";
    tmp(06592) := x"0000";
    tmp(06593) := x"0020";
    tmp(06594) := x"0820";
    tmp(06595) := x"0881";
    tmp(06596) := x"0880";
    tmp(06597) := x"0880";
    tmp(06598) := x"0880";
    tmp(06599) := x"0880";
    tmp(06600) := x"0880";
    tmp(06601) := x"0880";
    tmp(06602) := x"0040";
    tmp(06603) := x"0000";
    tmp(06604) := x"0000";
    tmp(06605) := x"0000";
    tmp(06606) := x"0000";
    tmp(06607) := x"0000";
    tmp(06608) := x"0000";
    tmp(06609) := x"0000";
    tmp(06610) := x"0000";
    tmp(06611) := x"0000";
    tmp(06612) := x"0000";
    tmp(06613) := x"0000";
    tmp(06614) := x"0000";
    tmp(06615) := x"0000";
    tmp(06616) := x"0020";
    tmp(06617) := x"0821";
    tmp(06618) := x"0841";
    tmp(06619) := x"0841";
    tmp(06620) := x"0821";
    tmp(06621) := x"0020";
    tmp(06622) := x"0841";
    tmp(06623) := x"0881";
    tmp(06624) := x"0880";
    tmp(06625) := x"0880";
    tmp(06626) := x"0880";
    tmp(06627) := x"0880";
    tmp(06628) := x"0880";
    tmp(06629) := x"0880";
    tmp(06630) := x"0860";
    tmp(06631) := x"0880";
    tmp(06632) := x"0860";
    tmp(06633) := x"0860";
    tmp(06634) := x"0880";
    tmp(06635) := x"0860";
    tmp(06636) := x"0860";
    tmp(06637) := x"0880";
    tmp(06638) := x"0880";
    tmp(06639) := x"0880";
    tmp(06640) := x"0880";
    tmp(06641) := x"0880";
    tmp(06642) := x"0880";
    tmp(06643) := x"0880";
    tmp(06644) := x"0880";
    tmp(06645) := x"0880";
    tmp(06646) := x"0880";
    tmp(06647) := x"08a0";
    tmp(06648) := x"08a0";
    tmp(06649) := x"08a0";
    tmp(06650) := x"08a0";
    tmp(06651) := x"08a0";
    tmp(06652) := x"08a0";
    tmp(06653) := x"08a0";
    tmp(06654) := x"08a0";
    tmp(06655) := x"08a0";
    tmp(06656) := x"08a0";
    tmp(06657) := x"08a0";
    tmp(06658) := x"08a0";
    tmp(06659) := x"08c0";
    tmp(06660) := x"08c0";
    tmp(06661) := x"08a0";
    tmp(06662) := x"08c0";
    tmp(06663) := x"08c0";
    tmp(06664) := x"08c0";
    tmp(06665) := x"08c0";
    tmp(06666) := x"08c0";
    tmp(06667) := x"08c0";
    tmp(06668) := x"08c0";
    tmp(06669) := x"08c0";
    tmp(06670) := x"08c0";
    tmp(06671) := x"08a0";
    tmp(06672) := x"08c0";
    tmp(06673) := x"08c0";
    tmp(06674) := x"08a0";
    tmp(06675) := x"08a0";
    tmp(06676) := x"08a0";
    tmp(06677) := x"ffff";
    tmp(06678) := x"ffff";
    tmp(06679) := x"ffff";
    tmp(06680) := x"ffff";
    tmp(06681) := x"ffff";
    tmp(06682) := x"ffff";
    tmp(06683) := x"ffff";
    tmp(06684) := x"ffff";
    tmp(06685) := x"ffff";
    tmp(06686) := x"ffff";
    tmp(06687) := x"ffff";
    tmp(06688) := x"ffff";
    tmp(06689) := x"ffff";
    tmp(06690) := x"ffff";
    tmp(06691) := x"ffff";
    tmp(06692) := x"ffff";
    tmp(06693) := x"ffff";
    tmp(06694) := x"ffff";
    tmp(06695) := x"ffff";
    tmp(06696) := x"ffff";
    tmp(06697) := x"ffff";
    tmp(06698) := x"ffff";
    tmp(06699) := x"ffff";
    tmp(06700) := x"ffff";
    tmp(06701) := x"ffff";
    tmp(06702) := x"ffff";
    tmp(06703) := x"ffff";
    tmp(06704) := x"ffff";
    tmp(06705) := x"ffff";
    tmp(06706) := x"ffff";
    tmp(06707) := x"ffff";
    tmp(06708) := x"ffff";
    tmp(06709) := x"ffff";
    tmp(06710) := x"ffff";
    tmp(06711) := x"ffff";
    tmp(06712) := x"ffff";
    tmp(06713) := x"ffff";
    tmp(06714) := x"ffff";
    tmp(06715) := x"ffff";
    tmp(06716) := x"ffff";
    tmp(06717) := x"0820";
    tmp(06718) := x"0820";
    tmp(06719) := x"0820";
    tmp(06720) := x"0000";
    tmp(06721) := x"0020";
    tmp(06722) := x"0020";
    tmp(06723) := x"0020";
    tmp(06724) := x"0020";
    tmp(06725) := x"0040";
    tmp(06726) := x"0040";
    tmp(06727) := x"0040";
    tmp(06728) := x"0040";
    tmp(06729) := x"0040";
    tmp(06730) := x"0040";
    tmp(06731) := x"0040";
    tmp(06732) := x"0040";
    tmp(06733) := x"0840";
    tmp(06734) := x"0840";
    tmp(06735) := x"0840";
    tmp(06736) := x"0840";
    tmp(06737) := x"0840";
    tmp(06738) := x"0840";
    tmp(06739) := x"0820";
    tmp(06740) := x"0820";
    tmp(06741) := x"0820";
    tmp(06742) := x"0820";
    tmp(06743) := x"0820";
    tmp(06744) := x"0820";
    tmp(06745) := x"0820";
    tmp(06746) := x"0820";
    tmp(06747) := x"0820";
    tmp(06748) := x"0820";
    tmp(06749) := x"0820";
    tmp(06750) := x"0820";
    tmp(06751) := x"0820";
    tmp(06752) := x"0820";
    tmp(06753) := x"0820";
    tmp(06754) := x"0820";
    tmp(06755) := x"0820";
    tmp(06756) := x"0820";
    tmp(06757) := x"0820";
    tmp(06758) := x"0820";
    tmp(06759) := x"0820";
    tmp(06760) := x"0820";
    tmp(06761) := x"0820";
    tmp(06762) := x"0820";
    tmp(06763) := x"0820";
    tmp(06764) := x"0840";
    tmp(06765) := x"0840";
    tmp(06766) := x"0840";
    tmp(06767) := x"0840";
    tmp(06768) := x"0840";
    tmp(06769) := x"0840";
    tmp(06770) := x"0840";
    tmp(06771) := x"0840";
    tmp(06772) := x"0840";
    tmp(06773) := x"0840";
    tmp(06774) := x"0840";
    tmp(06775) := x"0840";
    tmp(06776) := x"0840";
    tmp(06777) := x"0840";
    tmp(06778) := x"0840";
    tmp(06779) := x"0840";
    tmp(06780) := x"0841";
    tmp(06781) := x"0840";
    tmp(06782) := x"0840";
    tmp(06783) := x"0841";
    tmp(06784) := x"0840";
    tmp(06785) := x"0840";
    tmp(06786) := x"0840";
    tmp(06787) := x"0840";
    tmp(06788) := x"0840";
    tmp(06789) := x"0840";
    tmp(06790) := x"0840";
    tmp(06791) := x"0840";
    tmp(06792) := x"0840";
    tmp(06793) := x"0840";
    tmp(06794) := x"0840";
    tmp(06795) := x"0840";
    tmp(06796) := x"0840";
    tmp(06797) := x"0840";
    tmp(06798) := x"0840";
    tmp(06799) := x"0840";
    tmp(06800) := x"0840";
    tmp(06801) := x"0840";
    tmp(06802) := x"0840";
    tmp(06803) := x"0840";
    tmp(06804) := x"0840";
    tmp(06805) := x"0860";
    tmp(06806) := x"0860";
    tmp(06807) := x"0860";
    tmp(06808) := x"0860";
    tmp(06809) := x"0860";
    tmp(06810) := x"0860";
    tmp(06811) := x"0860";
    tmp(06812) := x"0860";
    tmp(06813) := x"0860";
    tmp(06814) := x"0880";
    tmp(06815) := x"0880";
    tmp(06816) := x"0880";
    tmp(06817) := x"0880";
    tmp(06818) := x"0880";
    tmp(06819) := x"0880";
    tmp(06820) := x"0880";
    tmp(06821) := x"08a0";
    tmp(06822) := x"08a0";
    tmp(06823) := x"08a0";
    tmp(06824) := x"08a0";
    tmp(06825) := x"0860";
    tmp(06826) := x"0020";
    tmp(06827) := x"0000";
    tmp(06828) := x"0000";
    tmp(06829) := x"0000";
    tmp(06830) := x"0000";
    tmp(06831) := x"0000";
    tmp(06832) := x"0020";
    tmp(06833) := x"0000";
    tmp(06834) := x"0000";
    tmp(06835) := x"0000";
    tmp(06836) := x"0020";
    tmp(06837) := x"0840";
    tmp(06838) := x"0880";
    tmp(06839) := x"0880";
    tmp(06840) := x"0880";
    tmp(06841) := x"0860";
    tmp(06842) := x"0020";
    tmp(06843) := x"0000";
    tmp(06844) := x"0000";
    tmp(06845) := x"0000";
    tmp(06846) := x"0000";
    tmp(06847) := x"0000";
    tmp(06848) := x"0000";
    tmp(06849) := x"0000";
    tmp(06850) := x"0000";
    tmp(06851) := x"0000";
    tmp(06852) := x"0000";
    tmp(06853) := x"0000";
    tmp(06854) := x"0000";
    tmp(06855) := x"0000";
    tmp(06856) := x"0020";
    tmp(06857) := x"0020";
    tmp(06858) := x"0821";
    tmp(06859) := x"0841";
    tmp(06860) := x"0841";
    tmp(06861) := x"0821";
    tmp(06862) := x"0020";
    tmp(06863) := x"0841";
    tmp(06864) := x"0880";
    tmp(06865) := x"0880";
    tmp(06866) := x"0880";
    tmp(06867) := x"0880";
    tmp(06868) := x"0880";
    tmp(06869) := x"0880";
    tmp(06870) := x"0860";
    tmp(06871) := x"0860";
    tmp(06872) := x"0860";
    tmp(06873) := x"0860";
    tmp(06874) := x"0860";
    tmp(06875) := x"0860";
    tmp(06876) := x"0860";
    tmp(06877) := x"0860";
    tmp(06878) := x"0860";
    tmp(06879) := x"0860";
    tmp(06880) := x"0860";
    tmp(06881) := x"0860";
    tmp(06882) := x"0860";
    tmp(06883) := x"0860";
    tmp(06884) := x"0860";
    tmp(06885) := x"0860";
    tmp(06886) := x"0880";
    tmp(06887) := x"0880";
    tmp(06888) := x"0880";
    tmp(06889) := x"0880";
    tmp(06890) := x"0880";
    tmp(06891) := x"0880";
    tmp(06892) := x"0880";
    tmp(06893) := x"0880";
    tmp(06894) := x"0880";
    tmp(06895) := x"08a0";
    tmp(06896) := x"08a0";
    tmp(06897) := x"08a0";
    tmp(06898) := x"08a0";
    tmp(06899) := x"08a0";
    tmp(06900) := x"08a0";
    tmp(06901) := x"08a0";
    tmp(06902) := x"08a0";
    tmp(06903) := x"08a0";
    tmp(06904) := x"08a0";
    tmp(06905) := x"08a0";
    tmp(06906) := x"08a0";
    tmp(06907) := x"08a0";
    tmp(06908) := x"08a0";
    tmp(06909) := x"08a0";
    tmp(06910) := x"08a0";
    tmp(06911) := x"08a0";
    tmp(06912) := x"08a0";
    tmp(06913) := x"08a0";
    tmp(06914) := x"08a0";
    tmp(06915) := x"08a0";
    tmp(06916) := x"08a0";
    tmp(06917) := x"ffff";
    tmp(06918) := x"ffff";
    tmp(06919) := x"ffff";
    tmp(06920) := x"ffff";
    tmp(06921) := x"ffff";
    tmp(06922) := x"ffff";
    tmp(06923) := x"ffff";
    tmp(06924) := x"ffff";
    tmp(06925) := x"ffff";
    tmp(06926) := x"ffff";
    tmp(06927) := x"ffff";
    tmp(06928) := x"ffff";
    tmp(06929) := x"ffff";
    tmp(06930) := x"ffff";
    tmp(06931) := x"ffff";
    tmp(06932) := x"ffff";
    tmp(06933) := x"ffff";
    tmp(06934) := x"ffff";
    tmp(06935) := x"ffff";
    tmp(06936) := x"ffff";
    tmp(06937) := x"ffff";
    tmp(06938) := x"ffff";
    tmp(06939) := x"ffff";
    tmp(06940) := x"ffff";
    tmp(06941) := x"ffff";
    tmp(06942) := x"ffff";
    tmp(06943) := x"ffff";
    tmp(06944) := x"ffff";
    tmp(06945) := x"ffff";
    tmp(06946) := x"ffff";
    tmp(06947) := x"ffff";
    tmp(06948) := x"ffff";
    tmp(06949) := x"ffff";
    tmp(06950) := x"ffff";
    tmp(06951) := x"ffff";
    tmp(06952) := x"ffff";
    tmp(06953) := x"ffff";
    tmp(06954) := x"ffff";
    tmp(06955) := x"ffff";
    tmp(06956) := x"ffff";
    tmp(06957) := x"0820";
    tmp(06958) := x"0820";
    tmp(06959) := x"0820";
    tmp(06960) := x"0000";
    tmp(06961) := x"0020";
    tmp(06962) := x"0020";
    tmp(06963) := x"0020";
    tmp(06964) := x"0040";
    tmp(06965) := x"0040";
    tmp(06966) := x"0040";
    tmp(06967) := x"0040";
    tmp(06968) := x"0040";
    tmp(06969) := x"0040";
    tmp(06970) := x"0040";
    tmp(06971) := x"0040";
    tmp(06972) := x"0840";
    tmp(06973) := x"0840";
    tmp(06974) := x"0840";
    tmp(06975) := x"0840";
    tmp(06976) := x"0840";
    tmp(06977) := x"0840";
    tmp(06978) := x"0820";
    tmp(06979) := x"0820";
    tmp(06980) := x"0820";
    tmp(06981) := x"0820";
    tmp(06982) := x"0820";
    tmp(06983) := x"0820";
    tmp(06984) := x"0820";
    tmp(06985) := x"0820";
    tmp(06986) := x"0820";
    tmp(06987) := x"0820";
    tmp(06988) := x"0820";
    tmp(06989) := x"0820";
    tmp(06990) := x"0820";
    tmp(06991) := x"0820";
    tmp(06992) := x"0820";
    tmp(06993) := x"0820";
    tmp(06994) := x"0820";
    tmp(06995) := x"0820";
    tmp(06996) := x"0820";
    tmp(06997) := x"0820";
    tmp(06998) := x"0820";
    tmp(06999) := x"0820";
    tmp(07000) := x"0820";
    tmp(07001) := x"0820";
    tmp(07002) := x"0840";
    tmp(07003) := x"0840";
    tmp(07004) := x"0840";
    tmp(07005) := x"0840";
    tmp(07006) := x"0840";
    tmp(07007) := x"0840";
    tmp(07008) := x"0840";
    tmp(07009) := x"0840";
    tmp(07010) := x"0840";
    tmp(07011) := x"0840";
    tmp(07012) := x"0840";
    tmp(07013) := x"0840";
    tmp(07014) := x"0840";
    tmp(07015) := x"0840";
    tmp(07016) := x"0840";
    tmp(07017) := x"0840";
    tmp(07018) := x"0840";
    tmp(07019) := x"0840";
    tmp(07020) := x"0840";
    tmp(07021) := x"0840";
    tmp(07022) := x"0840";
    tmp(07023) := x"0840";
    tmp(07024) := x"0840";
    tmp(07025) := x"0840";
    tmp(07026) := x"0840";
    tmp(07027) := x"0841";
    tmp(07028) := x"0841";
    tmp(07029) := x"0840";
    tmp(07030) := x"0840";
    tmp(07031) := x"0840";
    tmp(07032) := x"0840";
    tmp(07033) := x"0840";
    tmp(07034) := x"0840";
    tmp(07035) := x"0840";
    tmp(07036) := x"0840";
    tmp(07037) := x"0840";
    tmp(07038) := x"0840";
    tmp(07039) := x"0840";
    tmp(07040) := x"0840";
    tmp(07041) := x"0840";
    tmp(07042) := x"0840";
    tmp(07043) := x"0840";
    tmp(07044) := x"0860";
    tmp(07045) := x"0860";
    tmp(07046) := x"0860";
    tmp(07047) := x"0860";
    tmp(07048) := x"0860";
    tmp(07049) := x"0860";
    tmp(07050) := x"0860";
    tmp(07051) := x"0860";
    tmp(07052) := x"0860";
    tmp(07053) := x"0860";
    tmp(07054) := x"0880";
    tmp(07055) := x"0880";
    tmp(07056) := x"0880";
    tmp(07057) := x"0880";
    tmp(07058) := x"0880";
    tmp(07059) := x"0880";
    tmp(07060) := x"0880";
    tmp(07061) := x"0880";
    tmp(07062) := x"0880";
    tmp(07063) := x"0880";
    tmp(07064) := x"0860";
    tmp(07065) := x"0020";
    tmp(07066) := x"0000";
    tmp(07067) := x"0000";
    tmp(07068) := x"0000";
    tmp(07069) := x"0000";
    tmp(07070) := x"0000";
    tmp(07071) := x"0000";
    tmp(07072) := x"0020";
    tmp(07073) := x"0000";
    tmp(07074) := x"0000";
    tmp(07075) := x"0000";
    tmp(07076) := x"0000";
    tmp(07077) := x"0000";
    tmp(07078) := x"0020";
    tmp(07079) := x"0860";
    tmp(07080) := x"0880";
    tmp(07081) := x"0840";
    tmp(07082) := x"0000";
    tmp(07083) := x"0000";
    tmp(07084) := x"0000";
    tmp(07085) := x"0000";
    tmp(07086) := x"0000";
    tmp(07087) := x"0000";
    tmp(07088) := x"0000";
    tmp(07089) := x"0000";
    tmp(07090) := x"0000";
    tmp(07091) := x"0000";
    tmp(07092) := x"0000";
    tmp(07093) := x"0000";
    tmp(07094) := x"0000";
    tmp(07095) := x"0020";
    tmp(07096) := x"0000";
    tmp(07097) := x"0020";
    tmp(07098) := x"0021";
    tmp(07099) := x"0841";
    tmp(07100) := x"0841";
    tmp(07101) := x"0841";
    tmp(07102) := x"0821";
    tmp(07103) := x"0020";
    tmp(07104) := x"0861";
    tmp(07105) := x"0880";
    tmp(07106) := x"0880";
    tmp(07107) := x"0880";
    tmp(07108) := x"0880";
    tmp(07109) := x"0860";
    tmp(07110) := x"0880";
    tmp(07111) := x"0860";
    tmp(07112) := x"0860";
    tmp(07113) := x"0860";
    tmp(07114) := x"0860";
    tmp(07115) := x"0860";
    tmp(07116) := x"0860";
    tmp(07117) := x"0860";
    tmp(07118) := x"0860";
    tmp(07119) := x"0860";
    tmp(07120) := x"0860";
    tmp(07121) := x"0860";
    tmp(07122) := x"0860";
    tmp(07123) := x"0860";
    tmp(07124) := x"0860";
    tmp(07125) := x"0860";
    tmp(07126) := x"0860";
    tmp(07127) := x"0860";
    tmp(07128) := x"0860";
    tmp(07129) := x"0860";
    tmp(07130) := x"0860";
    tmp(07131) := x"0860";
    tmp(07132) := x"0860";
    tmp(07133) := x"0060";
    tmp(07134) := x"0060";
    tmp(07135) := x"0860";
    tmp(07136) := x"0060";
    tmp(07137) := x"0880";
    tmp(07138) := x"0880";
    tmp(07139) := x"0880";
    tmp(07140) := x"0880";
    tmp(07141) := x"0880";
    tmp(07142) := x"0880";
    tmp(07143) := x"0880";
    tmp(07144) := x"08a0";
    tmp(07145) := x"0880";
    tmp(07146) := x"08a0";
    tmp(07147) := x"08a0";
    tmp(07148) := x"08a0";
    tmp(07149) := x"08a0";
    tmp(07150) := x"08a0";
    tmp(07151) := x"08a0";
    tmp(07152) := x"00a0";
    tmp(07153) := x"08a0";
    tmp(07154) := x"08a0";
    tmp(07155) := x"08a0";
    tmp(07156) := x"00a0";
    tmp(07157) := x"ffff";
    tmp(07158) := x"ffff";
    tmp(07159) := x"ffff";
    tmp(07160) := x"ffff";
    tmp(07161) := x"ffff";
    tmp(07162) := x"ffff";
    tmp(07163) := x"ffff";
    tmp(07164) := x"ffff";
    tmp(07165) := x"ffff";
    tmp(07166) := x"ffff";
    tmp(07167) := x"ffff";
    tmp(07168) := x"ffff";
    tmp(07169) := x"ffff";
    tmp(07170) := x"ffff";
    tmp(07171) := x"ffff";
    tmp(07172) := x"ffff";
    tmp(07173) := x"ffff";
    tmp(07174) := x"ffff";
    tmp(07175) := x"ffff";
    tmp(07176) := x"ffff";
    tmp(07177) := x"ffff";
    tmp(07178) := x"ffff";
    tmp(07179) := x"ffff";
    tmp(07180) := x"ffff";
    tmp(07181) := x"ffff";
    tmp(07182) := x"ffff";
    tmp(07183) := x"ffff";
    tmp(07184) := x"ffff";
    tmp(07185) := x"ffff";
    tmp(07186) := x"ffff";
    tmp(07187) := x"ffff";
    tmp(07188) := x"ffff";
    tmp(07189) := x"ffff";
    tmp(07190) := x"ffff";
    tmp(07191) := x"ffff";
    tmp(07192) := x"ffff";
    tmp(07193) := x"ffff";
    tmp(07194) := x"ffff";
    tmp(07195) := x"ffff";
    tmp(07196) := x"ffff";
    tmp(07197) := x"0820";
    tmp(07198) := x"0820";
    tmp(07199) := x"0820";
    tmp(07200) := x"0000";
    tmp(07201) := x"0020";
    tmp(07202) := x"0020";
    tmp(07203) := x"0040";
    tmp(07204) := x"0040";
    tmp(07205) := x"0040";
    tmp(07206) := x"0040";
    tmp(07207) := x"0040";
    tmp(07208) := x"0040";
    tmp(07209) := x"0040";
    tmp(07210) := x"0040";
    tmp(07211) := x"0840";
    tmp(07212) := x"0840";
    tmp(07213) := x"0840";
    tmp(07214) := x"0840";
    tmp(07215) := x"0840";
    tmp(07216) := x"0820";
    tmp(07217) := x"0820";
    tmp(07218) := x"0820";
    tmp(07219) := x"0820";
    tmp(07220) := x"0820";
    tmp(07221) := x"0820";
    tmp(07222) := x"0820";
    tmp(07223) := x"0820";
    tmp(07224) := x"0820";
    tmp(07225) := x"0820";
    tmp(07226) := x"0820";
    tmp(07227) := x"0820";
    tmp(07228) := x"0820";
    tmp(07229) := x"0820";
    tmp(07230) := x"0820";
    tmp(07231) := x"0820";
    tmp(07232) := x"0820";
    tmp(07233) := x"0820";
    tmp(07234) := x"0820";
    tmp(07235) := x"0820";
    tmp(07236) := x"0820";
    tmp(07237) := x"0820";
    tmp(07238) := x"0820";
    tmp(07239) := x"0820";
    tmp(07240) := x"0820";
    tmp(07241) := x"0820";
    tmp(07242) := x"0840";
    tmp(07243) := x"0840";
    tmp(07244) := x"0840";
    tmp(07245) := x"0840";
    tmp(07246) := x"0840";
    tmp(07247) := x"0840";
    tmp(07248) := x"0840";
    tmp(07249) := x"0840";
    tmp(07250) := x"0840";
    tmp(07251) := x"0840";
    tmp(07252) := x"0840";
    tmp(07253) := x"0840";
    tmp(07254) := x"0840";
    tmp(07255) := x"0840";
    tmp(07256) := x"0840";
    tmp(07257) := x"0840";
    tmp(07258) := x"0841";
    tmp(07259) := x"0840";
    tmp(07260) := x"0841";
    tmp(07261) := x"0840";
    tmp(07262) := x"0841";
    tmp(07263) := x"0841";
    tmp(07264) := x"0840";
    tmp(07265) := x"0840";
    tmp(07266) := x"0840";
    tmp(07267) := x"0841";
    tmp(07268) := x"0840";
    tmp(07269) := x"0840";
    tmp(07270) := x"0841";
    tmp(07271) := x"0840";
    tmp(07272) := x"0840";
    tmp(07273) := x"0840";
    tmp(07274) := x"0840";
    tmp(07275) := x"0840";
    tmp(07276) := x"0840";
    tmp(07277) := x"0840";
    tmp(07278) := x"0840";
    tmp(07279) := x"0840";
    tmp(07280) := x"0840";
    tmp(07281) := x"0840";
    tmp(07282) := x"0840";
    tmp(07283) := x"0860";
    tmp(07284) := x"0860";
    tmp(07285) := x"0860";
    tmp(07286) := x"0860";
    tmp(07287) := x"0860";
    tmp(07288) := x"0860";
    tmp(07289) := x"0860";
    tmp(07290) := x"0860";
    tmp(07291) := x"0860";
    tmp(07292) := x"0860";
    tmp(07293) := x"0880";
    tmp(07294) := x"0880";
    tmp(07295) := x"0880";
    tmp(07296) := x"0880";
    tmp(07297) := x"0880";
    tmp(07298) := x"0880";
    tmp(07299) := x"0880";
    tmp(07300) := x"0880";
    tmp(07301) := x"0880";
    tmp(07302) := x"0880";
    tmp(07303) := x"0880";
    tmp(07304) := x"0020";
    tmp(07305) := x"0000";
    tmp(07306) := x"0000";
    tmp(07307) := x"0000";
    tmp(07308) := x"0000";
    tmp(07309) := x"0000";
    tmp(07310) := x"0000";
    tmp(07311) := x"0020";
    tmp(07312) := x"0000";
    tmp(07313) := x"0000";
    tmp(07314) := x"0000";
    tmp(07315) := x"0000";
    tmp(07316) := x"0000";
    tmp(07317) := x"0000";
    tmp(07318) := x"0000";
    tmp(07319) := x"0000";
    tmp(07320) := x"0840";
    tmp(07321) := x"0020";
    tmp(07322) := x"0000";
    tmp(07323) := x"0000";
    tmp(07324) := x"0000";
    tmp(07325) := x"0000";
    tmp(07326) := x"0000";
    tmp(07327) := x"0000";
    tmp(07328) := x"0000";
    tmp(07329) := x"0000";
    tmp(07330) := x"0000";
    tmp(07331) := x"0000";
    tmp(07332) := x"0000";
    tmp(07333) := x"0000";
    tmp(07334) := x"0000";
    tmp(07335) := x"0020";
    tmp(07336) := x"0020";
    tmp(07337) := x"0020";
    tmp(07338) := x"0020";
    tmp(07339) := x"0021";
    tmp(07340) := x"0841";
    tmp(07341) := x"0841";
    tmp(07342) := x"0841";
    tmp(07343) := x"0821";
    tmp(07344) := x"0820";
    tmp(07345) := x"0861";
    tmp(07346) := x"0880";
    tmp(07347) := x"0880";
    tmp(07348) := x"0880";
    tmp(07349) := x"0880";
    tmp(07350) := x"0880";
    tmp(07351) := x"0860";
    tmp(07352) := x"0880";
    tmp(07353) := x"0860";
    tmp(07354) := x"0860";
    tmp(07355) := x"0860";
    tmp(07356) := x"0860";
    tmp(07357) := x"0860";
    tmp(07358) := x"0860";
    tmp(07359) := x"0860";
    tmp(07360) := x"0860";
    tmp(07361) := x"0860";
    tmp(07362) := x"0860";
    tmp(07363) := x"0840";
    tmp(07364) := x"0860";
    tmp(07365) := x"0860";
    tmp(07366) := x"0860";
    tmp(07367) := x"0860";
    tmp(07368) := x"0860";
    tmp(07369) := x"0860";
    tmp(07370) := x"0860";
    tmp(07371) := x"0860";
    tmp(07372) := x"0860";
    tmp(07373) := x"0860";
    tmp(07374) := x"0860";
    tmp(07375) := x"0060";
    tmp(07376) := x"0060";
    tmp(07377) := x"0060";
    tmp(07378) := x"0060";
    tmp(07379) := x"0860";
    tmp(07380) := x"0860";
    tmp(07381) := x"0060";
    tmp(07382) := x"0080";
    tmp(07383) := x"0880";
    tmp(07384) := x"0880";
    tmp(07385) := x"0880";
    tmp(07386) := x"0880";
    tmp(07387) := x"0080";
    tmp(07388) := x"0080";
    tmp(07389) := x"0080";
    tmp(07390) := x"0080";
    tmp(07391) := x"0080";
    tmp(07392) := x"0080";
    tmp(07393) := x"0080";
    tmp(07394) := x"0080";
    tmp(07395) := x"0080";
    tmp(07396) := x"0080";
    tmp(07397) := x"ffff";
    tmp(07398) := x"ffff";
    tmp(07399) := x"ffff";
    tmp(07400) := x"ffff";
    tmp(07401) := x"ffff";
    tmp(07402) := x"ffff";
    tmp(07403) := x"ffff";
    tmp(07404) := x"ffff";
    tmp(07405) := x"ffff";
    tmp(07406) := x"ffff";
    tmp(07407) := x"ffff";
    tmp(07408) := x"ffff";
    tmp(07409) := x"ffff";
    tmp(07410) := x"ffff";
    tmp(07411) := x"ffff";
    tmp(07412) := x"ffff";
    tmp(07413) := x"ffff";
    tmp(07414) := x"ffff";
    tmp(07415) := x"ffff";
    tmp(07416) := x"ffff";
    tmp(07417) := x"ffff";
    tmp(07418) := x"ffff";
    tmp(07419) := x"ffff";
    tmp(07420) := x"ffff";
    tmp(07421) := x"ffff";
    tmp(07422) := x"ffff";
    tmp(07423) := x"ffff";
    tmp(07424) := x"ffff";
    tmp(07425) := x"ffff";
    tmp(07426) := x"ffff";
    tmp(07427) := x"ffff";
    tmp(07428) := x"ffff";
    tmp(07429) := x"ffff";
    tmp(07430) := x"ffff";
    tmp(07431) := x"ffff";
    tmp(07432) := x"ffff";
    tmp(07433) := x"ffff";
    tmp(07434) := x"ffff";
    tmp(07435) := x"ffff";
    tmp(07436) := x"ffff";
    tmp(07437) := x"0820";
    tmp(07438) := x"0820";
    tmp(07439) := x"0820";
    tmp(07440) := x"0000";
    tmp(07441) := x"0040";
    tmp(07442) := x"0040";
    tmp(07443) := x"0040";
    tmp(07444) := x"0040";
    tmp(07445) := x"0040";
    tmp(07446) := x"0040";
    tmp(07447) := x"0040";
    tmp(07448) := x"0040";
    tmp(07449) := x"0040";
    tmp(07450) := x"0040";
    tmp(07451) := x"0840";
    tmp(07452) := x"0840";
    tmp(07453) := x"0840";
    tmp(07454) := x"0840";
    tmp(07455) := x"0820";
    tmp(07456) := x"0820";
    tmp(07457) := x"0820";
    tmp(07458) := x"0820";
    tmp(07459) := x"0820";
    tmp(07460) := x"0820";
    tmp(07461) := x"0820";
    tmp(07462) := x"0820";
    tmp(07463) := x"0820";
    tmp(07464) := x"0820";
    tmp(07465) := x"0820";
    tmp(07466) := x"0820";
    tmp(07467) := x"0820";
    tmp(07468) := x"0820";
    tmp(07469) := x"0820";
    tmp(07470) := x"0820";
    tmp(07471) := x"0820";
    tmp(07472) := x"0820";
    tmp(07473) := x"0820";
    tmp(07474) := x"0820";
    tmp(07475) := x"0820";
    tmp(07476) := x"0820";
    tmp(07477) := x"0820";
    tmp(07478) := x"0820";
    tmp(07479) := x"0820";
    tmp(07480) := x"0820";
    tmp(07481) := x"0820";
    tmp(07482) := x"0820";
    tmp(07483) := x"0840";
    tmp(07484) := x"0840";
    tmp(07485) := x"0840";
    tmp(07486) := x"0840";
    tmp(07487) := x"0840";
    tmp(07488) := x"0840";
    tmp(07489) := x"0840";
    tmp(07490) := x"0840";
    tmp(07491) := x"0840";
    tmp(07492) := x"0840";
    tmp(07493) := x"0840";
    tmp(07494) := x"0840";
    tmp(07495) := x"0840";
    tmp(07496) := x"0840";
    tmp(07497) := x"0840";
    tmp(07498) := x"0840";
    tmp(07499) := x"0840";
    tmp(07500) := x"0840";
    tmp(07501) := x"0840";
    tmp(07502) := x"0841";
    tmp(07503) := x"0841";
    tmp(07504) := x"0840";
    tmp(07505) := x"0840";
    tmp(07506) := x"0841";
    tmp(07507) := x"0841";
    tmp(07508) := x"0841";
    tmp(07509) := x"0841";
    tmp(07510) := x"0840";
    tmp(07511) := x"0840";
    tmp(07512) := x"0840";
    tmp(07513) := x"0840";
    tmp(07514) := x"0840";
    tmp(07515) := x"0840";
    tmp(07516) := x"0840";
    tmp(07517) := x"0840";
    tmp(07518) := x"0840";
    tmp(07519) := x"0840";
    tmp(07520) := x"0840";
    tmp(07521) := x"0840";
    tmp(07522) := x"0840";
    tmp(07523) := x"0860";
    tmp(07524) := x"0860";
    tmp(07525) := x"0860";
    tmp(07526) := x"0860";
    tmp(07527) := x"0860";
    tmp(07528) := x"0860";
    tmp(07529) := x"0860";
    tmp(07530) := x"0860";
    tmp(07531) := x"0860";
    tmp(07532) := x"0860";
    tmp(07533) := x"0880";
    tmp(07534) := x"0880";
    tmp(07535) := x"0880";
    tmp(07536) := x"0880";
    tmp(07537) := x"0880";
    tmp(07538) := x"0880";
    tmp(07539) := x"0880";
    tmp(07540) := x"0880";
    tmp(07541) := x"0880";
    tmp(07542) := x"0880";
    tmp(07543) := x"0020";
    tmp(07544) := x"0020";
    tmp(07545) := x"0000";
    tmp(07546) := x"0000";
    tmp(07547) := x"0000";
    tmp(07548) := x"0000";
    tmp(07549) := x"0000";
    tmp(07550) := x"0000";
    tmp(07551) := x"0020";
    tmp(07552) := x"0000";
    tmp(07553) := x"0000";
    tmp(07554) := x"0000";
    tmp(07555) := x"0000";
    tmp(07556) := x"0000";
    tmp(07557) := x"0000";
    tmp(07558) := x"0000";
    tmp(07559) := x"0000";
    tmp(07560) := x"0000";
    tmp(07561) := x"0000";
    tmp(07562) := x"0000";
    tmp(07563) := x"0000";
    tmp(07564) := x"0000";
    tmp(07565) := x"0000";
    tmp(07566) := x"0000";
    tmp(07567) := x"0000";
    tmp(07568) := x"0000";
    tmp(07569) := x"0000";
    tmp(07570) := x"0000";
    tmp(07571) := x"0000";
    tmp(07572) := x"0000";
    tmp(07573) := x"0000";
    tmp(07574) := x"0020";
    tmp(07575) := x"0020";
    tmp(07576) := x"0020";
    tmp(07577) := x"0020";
    tmp(07578) := x"0020";
    tmp(07579) := x"0020";
    tmp(07580) := x"0821";
    tmp(07581) := x"0841";
    tmp(07582) := x"0841";
    tmp(07583) := x"0841";
    tmp(07584) := x"0821";
    tmp(07585) := x"0841";
    tmp(07586) := x"0881";
    tmp(07587) := x"0880";
    tmp(07588) := x"0880";
    tmp(07589) := x"0880";
    tmp(07590) := x"0880";
    tmp(07591) := x"0880";
    tmp(07592) := x"0880";
    tmp(07593) := x"0860";
    tmp(07594) := x"0860";
    tmp(07595) := x"0860";
    tmp(07596) := x"0860";
    tmp(07597) := x"0860";
    tmp(07598) := x"0860";
    tmp(07599) := x"0860";
    tmp(07600) := x"0860";
    tmp(07601) := x"0860";
    tmp(07602) := x"0860";
    tmp(07603) := x"0840";
    tmp(07604) := x"0840";
    tmp(07605) := x"0840";
    tmp(07606) := x"0840";
    tmp(07607) := x"0840";
    tmp(07608) := x"0840";
    tmp(07609) := x"0840";
    tmp(07610) := x"0840";
    tmp(07611) := x"0840";
    tmp(07612) := x"0040";
    tmp(07613) := x"0840";
    tmp(07614) := x"0840";
    tmp(07615) := x"0040";
    tmp(07616) := x"0860";
    tmp(07617) := x"0060";
    tmp(07618) := x"0860";
    tmp(07619) := x"0060";
    tmp(07620) := x"0060";
    tmp(07621) := x"0060";
    tmp(07622) := x"0060";
    tmp(07623) := x"0060";
    tmp(07624) := x"0060";
    tmp(07625) := x"0060";
    tmp(07626) := x"0060";
    tmp(07627) := x"0060";
    tmp(07628) := x"0060";
    tmp(07629) := x"0060";
    tmp(07630) := x"0060";
    tmp(07631) := x"0060";
    tmp(07632) := x"0060";
    tmp(07633) := x"0060";
    tmp(07634) := x"0060";
    tmp(07635) := x"0080";
    tmp(07636) := x"0080";
    tmp(07637) := x"ffff";
    tmp(07638) := x"ffff";
    tmp(07639) := x"ffff";
    tmp(07640) := x"ffff";
    tmp(07641) := x"ffff";
    tmp(07642) := x"ffff";
    tmp(07643) := x"ffff";
    tmp(07644) := x"ffff";
    tmp(07645) := x"ffff";
    tmp(07646) := x"ffff";
    tmp(07647) := x"ffff";
    tmp(07648) := x"ffff";
    tmp(07649) := x"ffff";
    tmp(07650) := x"ffff";
    tmp(07651) := x"ffff";
    tmp(07652) := x"ffff";
    tmp(07653) := x"ffff";
    tmp(07654) := x"ffff";
    tmp(07655) := x"ffff";
    tmp(07656) := x"ffff";
    tmp(07657) := x"ffff";
    tmp(07658) := x"ffff";
    tmp(07659) := x"ffff";
    tmp(07660) := x"ffff";
    tmp(07661) := x"ffff";
    tmp(07662) := x"ffff";
    tmp(07663) := x"ffff";
    tmp(07664) := x"ffff";
    tmp(07665) := x"ffff";
    tmp(07666) := x"ffff";
    tmp(07667) := x"ffff";
    tmp(07668) := x"ffff";
    tmp(07669) := x"ffff";
    tmp(07670) := x"ffff";
    tmp(07671) := x"ffff";
    tmp(07672) := x"ffff";
    tmp(07673) := x"ffff";
    tmp(07674) := x"ffff";
    tmp(07675) := x"ffff";
    tmp(07676) := x"ffff";
    tmp(07677) := x"0820";
    tmp(07678) := x"0820";
    tmp(07679) := x"0820";
    tmp(07680) := x"0000";
    tmp(07681) := x"0040";
    tmp(07682) := x"0040";
    tmp(07683) := x"0040";
    tmp(07684) := x"0040";
    tmp(07685) := x"0040";
    tmp(07686) := x"0040";
    tmp(07687) := x"0040";
    tmp(07688) := x"0040";
    tmp(07689) := x"0040";
    tmp(07690) := x"0040";
    tmp(07691) := x"0840";
    tmp(07692) := x"0840";
    tmp(07693) := x"0840";
    tmp(07694) := x"0820";
    tmp(07695) := x"0820";
    tmp(07696) := x"0820";
    tmp(07697) := x"0820";
    tmp(07698) := x"0820";
    tmp(07699) := x"0820";
    tmp(07700) := x"0820";
    tmp(07701) := x"0820";
    tmp(07702) := x"0820";
    tmp(07703) := x"0820";
    tmp(07704) := x"0820";
    tmp(07705) := x"0820";
    tmp(07706) := x"0820";
    tmp(07707) := x"0820";
    tmp(07708) := x"0820";
    tmp(07709) := x"0820";
    tmp(07710) := x"0820";
    tmp(07711) := x"0820";
    tmp(07712) := x"0820";
    tmp(07713) := x"0820";
    tmp(07714) := x"0820";
    tmp(07715) := x"0820";
    tmp(07716) := x"0820";
    tmp(07717) := x"0820";
    tmp(07718) := x"0820";
    tmp(07719) := x"0820";
    tmp(07720) := x"0820";
    tmp(07721) := x"0820";
    tmp(07722) := x"0820";
    tmp(07723) := x"0840";
    tmp(07724) := x"0840";
    tmp(07725) := x"0840";
    tmp(07726) := x"0840";
    tmp(07727) := x"0840";
    tmp(07728) := x"0840";
    tmp(07729) := x"0840";
    tmp(07730) := x"0840";
    tmp(07731) := x"0840";
    tmp(07732) := x"0840";
    tmp(07733) := x"0840";
    tmp(07734) := x"0840";
    tmp(07735) := x"0841";
    tmp(07736) := x"0840";
    tmp(07737) := x"0840";
    tmp(07738) := x"0840";
    tmp(07739) := x"0840";
    tmp(07740) := x"0840";
    tmp(07741) := x"0840";
    tmp(07742) := x"0840";
    tmp(07743) := x"0841";
    tmp(07744) := x"0841";
    tmp(07745) := x"0841";
    tmp(07746) := x"0840";
    tmp(07747) := x"0841";
    tmp(07748) := x"0840";
    tmp(07749) := x"0841";
    tmp(07750) := x"0840";
    tmp(07751) := x"0840";
    tmp(07752) := x"0840";
    tmp(07753) := x"0840";
    tmp(07754) := x"0840";
    tmp(07755) := x"0840";
    tmp(07756) := x"0840";
    tmp(07757) := x"0840";
    tmp(07758) := x"0840";
    tmp(07759) := x"0840";
    tmp(07760) := x"0840";
    tmp(07761) := x"0840";
    tmp(07762) := x"0840";
    tmp(07763) := x"0860";
    tmp(07764) := x"0860";
    tmp(07765) := x"0860";
    tmp(07766) := x"0860";
    tmp(07767) := x"0860";
    tmp(07768) := x"0860";
    tmp(07769) := x"0860";
    tmp(07770) := x"0860";
    tmp(07771) := x"0860";
    tmp(07772) := x"0880";
    tmp(07773) := x"0880";
    tmp(07774) := x"0880";
    tmp(07775) := x"0880";
    tmp(07776) := x"0880";
    tmp(07777) := x"0880";
    tmp(07778) := x"0880";
    tmp(07779) := x"0880";
    tmp(07780) := x"0880";
    tmp(07781) := x"0880";
    tmp(07782) := x"0840";
    tmp(07783) := x"0000";
    tmp(07784) := x"0020";
    tmp(07785) := x"0000";
    tmp(07786) := x"0000";
    tmp(07787) := x"0000";
    tmp(07788) := x"0000";
    tmp(07789) := x"0000";
    tmp(07790) := x"0000";
    tmp(07791) := x"0020";
    tmp(07792) := x"0000";
    tmp(07793) := x"0000";
    tmp(07794) := x"0000";
    tmp(07795) := x"0000";
    tmp(07796) := x"0000";
    tmp(07797) := x"0000";
    tmp(07798) := x"0000";
    tmp(07799) := x"0000";
    tmp(07800) := x"0000";
    tmp(07801) := x"0000";
    tmp(07802) := x"0000";
    tmp(07803) := x"0000";
    tmp(07804) := x"0000";
    tmp(07805) := x"0000";
    tmp(07806) := x"0000";
    tmp(07807) := x"0000";
    tmp(07808) := x"0000";
    tmp(07809) := x"0000";
    tmp(07810) := x"0000";
    tmp(07811) := x"0020";
    tmp(07812) := x"0020";
    tmp(07813) := x"0000";
    tmp(07814) := x"0000";
    tmp(07815) := x"0020";
    tmp(07816) := x"0020";
    tmp(07817) := x"0020";
    tmp(07818) := x"0020";
    tmp(07819) := x"0020";
    tmp(07820) := x"0821";
    tmp(07821) := x"0841";
    tmp(07822) := x"0861";
    tmp(07823) := x"0861";
    tmp(07824) := x"0841";
    tmp(07825) := x"0820";
    tmp(07826) := x"0861";
    tmp(07827) := x"0880";
    tmp(07828) := x"0880";
    tmp(07829) := x"0880";
    tmp(07830) := x"0880";
    tmp(07831) := x"0880";
    tmp(07832) := x"0880";
    tmp(07833) := x"0860";
    tmp(07834) := x"0880";
    tmp(07835) := x"0860";
    tmp(07836) := x"0860";
    tmp(07837) := x"0860";
    tmp(07838) := x"0860";
    tmp(07839) := x"0860";
    tmp(07840) := x"0860";
    tmp(07841) := x"0860";
    tmp(07842) := x"0840";
    tmp(07843) := x"0840";
    tmp(07844) := x"0840";
    tmp(07845) := x"0840";
    tmp(07846) := x"0840";
    tmp(07847) := x"0840";
    tmp(07848) := x"0840";
    tmp(07849) := x"0840";
    tmp(07850) := x"0840";
    tmp(07851) := x"0840";
    tmp(07852) := x"0840";
    tmp(07853) := x"0040";
    tmp(07854) := x"0040";
    tmp(07855) := x"0040";
    tmp(07856) := x"0040";
    tmp(07857) := x"0040";
    tmp(07858) := x"0040";
    tmp(07859) := x"0040";
    tmp(07860) := x"0040";
    tmp(07861) := x"0040";
    tmp(07862) := x"0040";
    tmp(07863) := x"0040";
    tmp(07864) := x"0040";
    tmp(07865) := x"0040";
    tmp(07866) := x"0040";
    tmp(07867) := x"0040";
    tmp(07868) := x"0040";
    tmp(07869) := x"0040";
    tmp(07870) := x"0040";
    tmp(07871) := x"0040";
    tmp(07872) := x"0040";
    tmp(07873) := x"0040";
    tmp(07874) := x"0040";
    tmp(07875) := x"0060";
    tmp(07876) := x"0060";
    tmp(07877) := x"ffff";
    tmp(07878) := x"ffff";
    tmp(07879) := x"ffff";
    tmp(07880) := x"ffff";
    tmp(07881) := x"ffff";
    tmp(07882) := x"ffff";
    tmp(07883) := x"ffff";
    tmp(07884) := x"ffff";
    tmp(07885) := x"ffff";
    tmp(07886) := x"ffff";
    tmp(07887) := x"ffff";
    tmp(07888) := x"ffff";
    tmp(07889) := x"ffff";
    tmp(07890) := x"ffff";
    tmp(07891) := x"ffff";
    tmp(07892) := x"ffff";
    tmp(07893) := x"ffff";
    tmp(07894) := x"ffff";
    tmp(07895) := x"ffff";
    tmp(07896) := x"ffff";
    tmp(07897) := x"ffff";
    tmp(07898) := x"ffff";
    tmp(07899) := x"ffff";
    tmp(07900) := x"ffff";
    tmp(07901) := x"ffff";
    tmp(07902) := x"ffff";
    tmp(07903) := x"ffff";
    tmp(07904) := x"ffff";
    tmp(07905) := x"ffff";
    tmp(07906) := x"ffff";
    tmp(07907) := x"ffff";
    tmp(07908) := x"ffff";
    tmp(07909) := x"ffff";
    tmp(07910) := x"ffff";
    tmp(07911) := x"ffff";
    tmp(07912) := x"ffff";
    tmp(07913) := x"ffff";
    tmp(07914) := x"ffff";
    tmp(07915) := x"ffff";
    tmp(07916) := x"ffff";
    tmp(07917) := x"0820";
    tmp(07918) := x"0820";
    tmp(07919) := x"0820";
    tmp(07920) := x"0000";
    tmp(07921) := x"0040";
    tmp(07922) := x"0040";
    tmp(07923) := x"0040";
    tmp(07924) := x"0040";
    tmp(07925) := x"0040";
    tmp(07926) := x"0040";
    tmp(07927) := x"0040";
    tmp(07928) := x"0040";
    tmp(07929) := x"0040";
    tmp(07930) := x"0040";
    tmp(07931) := x"0840";
    tmp(07932) := x"0820";
    tmp(07933) := x"0020";
    tmp(07934) := x"0820";
    tmp(07935) := x"0820";
    tmp(07936) := x"0820";
    tmp(07937) := x"0820";
    tmp(07938) := x"0820";
    tmp(07939) := x"0820";
    tmp(07940) := x"0820";
    tmp(07941) := x"0820";
    tmp(07942) := x"0820";
    tmp(07943) := x"0820";
    tmp(07944) := x"0820";
    tmp(07945) := x"0820";
    tmp(07946) := x"0820";
    tmp(07947) := x"0820";
    tmp(07948) := x"0820";
    tmp(07949) := x"0820";
    tmp(07950) := x"0820";
    tmp(07951) := x"0820";
    tmp(07952) := x"0820";
    tmp(07953) := x"0820";
    tmp(07954) := x"0820";
    tmp(07955) := x"0820";
    tmp(07956) := x"0820";
    tmp(07957) := x"0820";
    tmp(07958) := x"0820";
    tmp(07959) := x"0820";
    tmp(07960) := x"0820";
    tmp(07961) := x"0820";
    tmp(07962) := x"0820";
    tmp(07963) := x"0840";
    tmp(07964) := x"0840";
    tmp(07965) := x"0840";
    tmp(07966) := x"0840";
    tmp(07967) := x"0840";
    tmp(07968) := x"0840";
    tmp(07969) := x"0840";
    tmp(07970) := x"0840";
    tmp(07971) := x"0840";
    tmp(07972) := x"0840";
    tmp(07973) := x"0840";
    tmp(07974) := x"0840";
    tmp(07975) := x"0840";
    tmp(07976) := x"0840";
    tmp(07977) := x"0840";
    tmp(07978) := x"0841";
    tmp(07979) := x"0841";
    tmp(07980) := x"0840";
    tmp(07981) := x"0840";
    tmp(07982) := x"0840";
    tmp(07983) := x"0840";
    tmp(07984) := x"0841";
    tmp(07985) := x"0841";
    tmp(07986) := x"0840";
    tmp(07987) := x"0840";
    tmp(07988) := x"0840";
    tmp(07989) := x"0840";
    tmp(07990) := x"0840";
    tmp(07991) := x"0840";
    tmp(07992) := x"0840";
    tmp(07993) := x"0840";
    tmp(07994) := x"0840";
    tmp(07995) := x"0840";
    tmp(07996) := x"0840";
    tmp(07997) := x"0840";
    tmp(07998) := x"0840";
    tmp(07999) := x"0840";
    tmp(08000) := x"0840";
    tmp(08001) := x"0840";
    tmp(08002) := x"0860";
    tmp(08003) := x"0860";
    tmp(08004) := x"0860";
    tmp(08005) := x"0860";
    tmp(08006) := x"0860";
    tmp(08007) := x"0860";
    tmp(08008) := x"0860";
    tmp(08009) := x"0860";
    tmp(08010) := x"0860";
    tmp(08011) := x"0860";
    tmp(08012) := x"0880";
    tmp(08013) := x"0880";
    tmp(08014) := x"0880";
    tmp(08015) := x"0880";
    tmp(08016) := x"0880";
    tmp(08017) := x"0880";
    tmp(08018) := x"0880";
    tmp(08019) := x"0880";
    tmp(08020) := x"0880";
    tmp(08021) := x"0880";
    tmp(08022) := x"0020";
    tmp(08023) := x"0000";
    tmp(08024) := x"0000";
    tmp(08025) := x"0000";
    tmp(08026) := x"0000";
    tmp(08027) := x"0000";
    tmp(08028) := x"0000";
    tmp(08029) := x"0000";
    tmp(08030) := x"0000";
    tmp(08031) := x"0020";
    tmp(08032) := x"0000";
    tmp(08033) := x"0000";
    tmp(08034) := x"0000";
    tmp(08035) := x"0000";
    tmp(08036) := x"0000";
    tmp(08037) := x"0000";
    tmp(08038) := x"0000";
    tmp(08039) := x"0000";
    tmp(08040) := x"0000";
    tmp(08041) := x"0000";
    tmp(08042) := x"0000";
    tmp(08043) := x"0000";
    tmp(08044) := x"0000";
    tmp(08045) := x"0000";
    tmp(08046) := x"0000";
    tmp(08047) := x"0000";
    tmp(08048) := x"0000";
    tmp(08049) := x"0000";
    tmp(08050) := x"0000";
    tmp(08051) := x"0000";
    tmp(08052) := x"0000";
    tmp(08053) := x"0000";
    tmp(08054) := x"0000";
    tmp(08055) := x"0000";
    tmp(08056) := x"0020";
    tmp(08057) := x"0020";
    tmp(08058) := x"0020";
    tmp(08059) := x"0020";
    tmp(08060) := x"0020";
    tmp(08061) := x"0821";
    tmp(08062) := x"0841";
    tmp(08063) := x"0861";
    tmp(08064) := x"0861";
    tmp(08065) := x"0861";
    tmp(08066) := x"0841";
    tmp(08067) := x"0881";
    tmp(08068) := x"0880";
    tmp(08069) := x"0880";
    tmp(08070) := x"0880";
    tmp(08071) := x"0880";
    tmp(08072) := x"0880";
    tmp(08073) := x"0880";
    tmp(08074) := x"0880";
    tmp(08075) := x"0880";
    tmp(08076) := x"0860";
    tmp(08077) := x"0860";
    tmp(08078) := x"0860";
    tmp(08079) := x"0860";
    tmp(08080) := x"0860";
    tmp(08081) := x"0860";
    tmp(08082) := x"0860";
    tmp(08083) := x"0860";
    tmp(08084) := x"0860";
    tmp(08085) := x"0840";
    tmp(08086) := x"0840";
    tmp(08087) := x"0840";
    tmp(08088) := x"0840";
    tmp(08089) := x"0840";
    tmp(08090) := x"0040";
    tmp(08091) := x"0840";
    tmp(08092) := x"0040";
    tmp(08093) := x"0040";
    tmp(08094) := x"0040";
    tmp(08095) := x"0040";
    tmp(08096) := x"0040";
    tmp(08097) := x"0040";
    tmp(08098) := x"0040";
    tmp(08099) := x"0040";
    tmp(08100) := x"0040";
    tmp(08101) := x"0040";
    tmp(08102) := x"0040";
    tmp(08103) := x"0040";
    tmp(08104) := x"0040";
    tmp(08105) := x"0040";
    tmp(08106) := x"0040";
    tmp(08107) := x"0040";
    tmp(08108) := x"0040";
    tmp(08109) := x"0040";
    tmp(08110) := x"0040";
    tmp(08111) := x"0040";
    tmp(08112) := x"0040";
    tmp(08113) := x"0040";
    tmp(08114) := x"0040";
    tmp(08115) := x"0040";
    tmp(08116) := x"0040";
    tmp(08117) := x"ffff";
    tmp(08118) := x"ffff";
    tmp(08119) := x"ffff";
    tmp(08120) := x"ffff";
    tmp(08121) := x"ffff";
    tmp(08122) := x"ffff";
    tmp(08123) := x"ffff";
    tmp(08124) := x"ffff";
    tmp(08125) := x"ffff";
    tmp(08126) := x"ffff";
    tmp(08127) := x"ffff";
    tmp(08128) := x"ffff";
    tmp(08129) := x"ffff";
    tmp(08130) := x"ffff";
    tmp(08131) := x"ffff";
    tmp(08132) := x"ffff";
    tmp(08133) := x"ffff";
    tmp(08134) := x"ffff";
    tmp(08135) := x"ffff";
    tmp(08136) := x"ffff";
    tmp(08137) := x"ffff";
    tmp(08138) := x"ffff";
    tmp(08139) := x"ffff";
    tmp(08140) := x"ffff";
    tmp(08141) := x"ffff";
    tmp(08142) := x"ffff";
    tmp(08143) := x"ffff";
    tmp(08144) := x"ffff";
    tmp(08145) := x"ffff";
    tmp(08146) := x"ffff";
    tmp(08147) := x"ffff";
    tmp(08148) := x"ffff";
    tmp(08149) := x"ffff";
    tmp(08150) := x"ffff";
    tmp(08151) := x"ffff";
    tmp(08152) := x"ffff";
    tmp(08153) := x"ffff";
    tmp(08154) := x"ffff";
    tmp(08155) := x"ffff";
    tmp(08156) := x"ffff";
    tmp(08157) := x"0820";
    tmp(08158) := x"0820";
    tmp(08159) := x"0820";
    tmp(08160) := x"0000";
    tmp(08161) := x"0040";
    tmp(08162) := x"0040";
    tmp(08163) := x"0040";
    tmp(08164) := x"0040";
    tmp(08165) := x"0040";
    tmp(08166) := x"0040";
    tmp(08167) := x"0040";
    tmp(08168) := x"0040";
    tmp(08169) := x"0040";
    tmp(08170) := x"0040";
    tmp(08171) := x"0840";
    tmp(08172) := x"0020";
    tmp(08173) := x"0020";
    tmp(08174) := x"0020";
    tmp(08175) := x"0020";
    tmp(08176) := x"0020";
    tmp(08177) := x"0020";
    tmp(08178) := x"0820";
    tmp(08179) := x"0020";
    tmp(08180) := x"0820";
    tmp(08181) := x"0820";
    tmp(08182) := x"0820";
    tmp(08183) := x"0820";
    tmp(08184) := x"0820";
    tmp(08185) := x"0820";
    tmp(08186) := x"0820";
    tmp(08187) := x"0820";
    tmp(08188) := x"0820";
    tmp(08189) := x"0820";
    tmp(08190) := x"0820";
    tmp(08191) := x"0820";
    tmp(08192) := x"0820";
    tmp(08193) := x"0820";
    tmp(08194) := x"0820";
    tmp(08195) := x"0820";
    tmp(08196) := x"0820";
    tmp(08197) := x"0820";
    tmp(08198) := x"0820";
    tmp(08199) := x"0820";
    tmp(08200) := x"0820";
    tmp(08201) := x"0820";
    tmp(08202) := x"0820";
    tmp(08203) := x"0820";
    tmp(08204) := x"0840";
    tmp(08205) := x"0840";
    tmp(08206) := x"0840";
    tmp(08207) := x"0840";
    tmp(08208) := x"0840";
    tmp(08209) := x"0840";
    tmp(08210) := x"0840";
    tmp(08211) := x"0840";
    tmp(08212) := x"0840";
    tmp(08213) := x"0840";
    tmp(08214) := x"0840";
    tmp(08215) := x"0840";
    tmp(08216) := x"0840";
    tmp(08217) := x"0840";
    tmp(08218) := x"0840";
    tmp(08219) := x"0841";
    tmp(08220) := x"0841";
    tmp(08221) := x"0841";
    tmp(08222) := x"0840";
    tmp(08223) := x"0841";
    tmp(08224) := x"0840";
    tmp(08225) := x"0840";
    tmp(08226) := x"0840";
    tmp(08227) := x"0841";
    tmp(08228) := x"0841";
    tmp(08229) := x"0841";
    tmp(08230) := x"0841";
    tmp(08231) := x"0841";
    tmp(08232) := x"0840";
    tmp(08233) := x"0840";
    tmp(08234) := x"0840";
    tmp(08235) := x"0840";
    tmp(08236) := x"0840";
    tmp(08237) := x"0840";
    tmp(08238) := x"0840";
    tmp(08239) := x"0840";
    tmp(08240) := x"0840";
    tmp(08241) := x"0840";
    tmp(08242) := x"0860";
    tmp(08243) := x"0860";
    tmp(08244) := x"0860";
    tmp(08245) := x"0860";
    tmp(08246) := x"0860";
    tmp(08247) := x"0860";
    tmp(08248) := x"0860";
    tmp(08249) := x"0860";
    tmp(08250) := x"0860";
    tmp(08251) := x"0880";
    tmp(08252) := x"0880";
    tmp(08253) := x"0880";
    tmp(08254) := x"0880";
    tmp(08255) := x"0880";
    tmp(08256) := x"0880";
    tmp(08257) := x"0880";
    tmp(08258) := x"0880";
    tmp(08259) := x"0880";
    tmp(08260) := x"0880";
    tmp(08261) := x"0860";
    tmp(08262) := x"0000";
    tmp(08263) := x"0000";
    tmp(08264) := x"0000";
    tmp(08265) := x"0000";
    tmp(08266) := x"0000";
    tmp(08267) := x"0000";
    tmp(08268) := x"0000";
    tmp(08269) := x"0000";
    tmp(08270) := x"0000";
    tmp(08271) := x"0820";
    tmp(08272) := x"0000";
    tmp(08273) := x"0000";
    tmp(08274) := x"0000";
    tmp(08275) := x"0000";
    tmp(08276) := x"0000";
    tmp(08277) := x"0000";
    tmp(08278) := x"0000";
    tmp(08279) := x"0020";
    tmp(08280) := x"0841";
    tmp(08281) := x"0821";
    tmp(08282) := x"0000";
    tmp(08283) := x"0000";
    tmp(08284) := x"0000";
    tmp(08285) := x"0000";
    tmp(08286) := x"0000";
    tmp(08287) := x"0000";
    tmp(08288) := x"0000";
    tmp(08289) := x"0000";
    tmp(08290) := x"0000";
    tmp(08291) := x"0000";
    tmp(08292) := x"0000";
    tmp(08293) := x"0000";
    tmp(08294) := x"0020";
    tmp(08295) := x"0020";
    tmp(08296) := x"0020";
    tmp(08297) := x"0020";
    tmp(08298) := x"0821";
    tmp(08299) := x"0020";
    tmp(08300) := x"0020";
    tmp(08301) := x"0020";
    tmp(08302) := x"0821";
    tmp(08303) := x"0841";
    tmp(08304) := x"0861";
    tmp(08305) := x"1081";
    tmp(08306) := x"1061";
    tmp(08307) := x"0861";
    tmp(08308) := x"08a0";
    tmp(08309) := x"08a0";
    tmp(08310) := x"08a0";
    tmp(08311) := x"0880";
    tmp(08312) := x"0880";
    tmp(08313) := x"0880";
    tmp(08314) := x"0880";
    tmp(08315) := x"0880";
    tmp(08316) := x"0880";
    tmp(08317) := x"0880";
    tmp(08318) := x"0880";
    tmp(08319) := x"0860";
    tmp(08320) := x"0860";
    tmp(08321) := x"0860";
    tmp(08322) := x"0860";
    tmp(08323) := x"0860";
    tmp(08324) := x"0860";
    tmp(08325) := x"0840";
    tmp(08326) := x"0840";
    tmp(08327) := x"0840";
    tmp(08328) := x"0840";
    tmp(08329) := x"0840";
    tmp(08330) := x"0840";
    tmp(08331) := x"0840";
    tmp(08332) := x"0840";
    tmp(08333) := x"0040";
    tmp(08334) := x"0020";
    tmp(08335) := x"0020";
    tmp(08336) := x"0020";
    tmp(08337) := x"0020";
    tmp(08338) := x"0020";
    tmp(08339) := x"0020";
    tmp(08340) := x"0020";
    tmp(08341) := x"0020";
    tmp(08342) := x"0020";
    tmp(08343) := x"0020";
    tmp(08344) := x"0020";
    tmp(08345) := x"0020";
    tmp(08346) := x"0020";
    tmp(08347) := x"0020";
    tmp(08348) := x"0020";
    tmp(08349) := x"0020";
    tmp(08350) := x"0020";
    tmp(08351) := x"0020";
    tmp(08352) := x"0020";
    tmp(08353) := x"0040";
    tmp(08354) := x"0020";
    tmp(08355) := x"0040";
    tmp(08356) := x"0020";
    tmp(08357) := x"ffff";
    tmp(08358) := x"ffff";
    tmp(08359) := x"ffff";
    tmp(08360) := x"ffff";
    tmp(08361) := x"ffff";
    tmp(08362) := x"ffff";
    tmp(08363) := x"ffff";
    tmp(08364) := x"ffff";
    tmp(08365) := x"ffff";
    tmp(08366) := x"ffff";
    tmp(08367) := x"ffff";
    tmp(08368) := x"ffff";
    tmp(08369) := x"ffff";
    tmp(08370) := x"ffff";
    tmp(08371) := x"ffff";
    tmp(08372) := x"ffff";
    tmp(08373) := x"ffff";
    tmp(08374) := x"ffff";
    tmp(08375) := x"ffff";
    tmp(08376) := x"ffff";
    tmp(08377) := x"ffff";
    tmp(08378) := x"ffff";
    tmp(08379) := x"ffff";
    tmp(08380) := x"ffff";
    tmp(08381) := x"ffff";
    tmp(08382) := x"ffff";
    tmp(08383) := x"ffff";
    tmp(08384) := x"ffff";
    tmp(08385) := x"ffff";
    tmp(08386) := x"ffff";
    tmp(08387) := x"ffff";
    tmp(08388) := x"ffff";
    tmp(08389) := x"ffff";
    tmp(08390) := x"ffff";
    tmp(08391) := x"ffff";
    tmp(08392) := x"ffff";
    tmp(08393) := x"ffff";
    tmp(08394) := x"ffff";
    tmp(08395) := x"ffff";
    tmp(08396) := x"ffff";
    tmp(08397) := x"0820";
    tmp(08398) := x"0820";
    tmp(08399) := x"0820";
    tmp(08400) := x"0000";
    tmp(08401) := x"0040";
    tmp(08402) := x"0040";
    tmp(08403) := x"0040";
    tmp(08404) := x"0040";
    tmp(08405) := x"0040";
    tmp(08406) := x"0040";
    tmp(08407) := x"0040";
    tmp(08408) := x"0040";
    tmp(08409) := x"0040";
    tmp(08410) := x"0040";
    tmp(08411) := x"0020";
    tmp(08412) := x"0020";
    tmp(08413) := x"0020";
    tmp(08414) := x"0020";
    tmp(08415) := x"0020";
    tmp(08416) := x"0020";
    tmp(08417) := x"0020";
    tmp(08418) := x"0020";
    tmp(08419) := x"0020";
    tmp(08420) := x"0020";
    tmp(08421) := x"0020";
    tmp(08422) := x"0820";
    tmp(08423) := x"0820";
    tmp(08424) := x"0820";
    tmp(08425) := x"0820";
    tmp(08426) := x"0820";
    tmp(08427) := x"0820";
    tmp(08428) := x"0820";
    tmp(08429) := x"0820";
    tmp(08430) := x"0820";
    tmp(08431) := x"0820";
    tmp(08432) := x"0820";
    tmp(08433) := x"0820";
    tmp(08434) := x"0820";
    tmp(08435) := x"0820";
    tmp(08436) := x"0820";
    tmp(08437) := x"0820";
    tmp(08438) := x"0820";
    tmp(08439) := x"0820";
    tmp(08440) := x"0820";
    tmp(08441) := x"0820";
    tmp(08442) := x"0840";
    tmp(08443) := x"0840";
    tmp(08444) := x"0840";
    tmp(08445) := x"0840";
    tmp(08446) := x"0840";
    tmp(08447) := x"0840";
    tmp(08448) := x"0840";
    tmp(08449) := x"0840";
    tmp(08450) := x"0840";
    tmp(08451) := x"0840";
    tmp(08452) := x"0840";
    tmp(08453) := x"0840";
    tmp(08454) := x"0840";
    tmp(08455) := x"0840";
    tmp(08456) := x"0840";
    tmp(08457) := x"0840";
    tmp(08458) := x"0840";
    tmp(08459) := x"0840";
    tmp(08460) := x"0840";
    tmp(08461) := x"0840";
    tmp(08462) := x"0840";
    tmp(08463) := x"0840";
    tmp(08464) := x"0840";
    tmp(08465) := x"0840";
    tmp(08466) := x"0840";
    tmp(08467) := x"0841";
    tmp(08468) := x"0841";
    tmp(08469) := x"0841";
    tmp(08470) := x"0840";
    tmp(08471) := x"0840";
    tmp(08472) := x"0840";
    tmp(08473) := x"0840";
    tmp(08474) := x"0840";
    tmp(08475) := x"0840";
    tmp(08476) := x"0840";
    tmp(08477) := x"0840";
    tmp(08478) := x"0840";
    tmp(08479) := x"0840";
    tmp(08480) := x"0840";
    tmp(08481) := x"0860";
    tmp(08482) := x"0860";
    tmp(08483) := x"0860";
    tmp(08484) := x"0860";
    tmp(08485) := x"0860";
    tmp(08486) := x"0860";
    tmp(08487) := x"0860";
    tmp(08488) := x"0860";
    tmp(08489) := x"0860";
    tmp(08490) := x"0880";
    tmp(08491) := x"0880";
    tmp(08492) := x"0880";
    tmp(08493) := x"0880";
    tmp(08494) := x"0880";
    tmp(08495) := x"0880";
    tmp(08496) := x"0880";
    tmp(08497) := x"0880";
    tmp(08498) := x"0880";
    tmp(08499) := x"0880";
    tmp(08500) := x"0880";
    tmp(08501) := x"0020";
    tmp(08502) := x"0000";
    tmp(08503) := x"0000";
    tmp(08504) := x"0000";
    tmp(08505) := x"0000";
    tmp(08506) := x"0000";
    tmp(08507) := x"0000";
    tmp(08508) := x"0000";
    tmp(08509) := x"0000";
    tmp(08510) := x"0000";
    tmp(08511) := x"0020";
    tmp(08512) := x"0021";
    tmp(08513) := x"0000";
    tmp(08514) := x"0000";
    tmp(08515) := x"0000";
    tmp(08516) := x"0000";
    tmp(08517) := x"0000";
    tmp(08518) := x"0000";
    tmp(08519) := x"0820";
    tmp(08520) := x"0020";
    tmp(08521) := x"0000";
    tmp(08522) := x"0000";
    tmp(08523) := x"0000";
    tmp(08524) := x"0000";
    tmp(08525) := x"0000";
    tmp(08526) := x"0000";
    tmp(08527) := x"0000";
    tmp(08528) := x"0000";
    tmp(08529) := x"0020";
    tmp(08530) := x"0000";
    tmp(08531) := x"0000";
    tmp(08532) := x"0020";
    tmp(08533) := x"0000";
    tmp(08534) := x"0000";
    tmp(08535) := x"0020";
    tmp(08536) := x"0020";
    tmp(08537) := x"0020";
    tmp(08538) := x"0821";
    tmp(08539) := x"0821";
    tmp(08540) := x"0821";
    tmp(08541) := x"0020";
    tmp(08542) := x"0020";
    tmp(08543) := x"0821";
    tmp(08544) := x"0841";
    tmp(08545) := x"1081";
    tmp(08546) := x"10a1";
    tmp(08547) := x"1061";
    tmp(08548) := x"10a1";
    tmp(08549) := x"08a0";
    tmp(08550) := x"08a0";
    tmp(08551) := x"08a0";
    tmp(08552) := x"08a0";
    tmp(08553) := x"08a0";
    tmp(08554) := x"08a0";
    tmp(08555) := x"08a0";
    tmp(08556) := x"0880";
    tmp(08557) := x"0880";
    tmp(08558) := x"0880";
    tmp(08559) := x"0880";
    tmp(08560) := x"0880";
    tmp(08561) := x"0880";
    tmp(08562) := x"0860";
    tmp(08563) := x"0860";
    tmp(08564) := x"0860";
    tmp(08565) := x"0860";
    tmp(08566) := x"0860";
    tmp(08567) := x"0860";
    tmp(08568) := x"0840";
    tmp(08569) := x"0840";
    tmp(08570) := x"0840";
    tmp(08571) := x"0840";
    tmp(08572) := x"0840";
    tmp(08573) := x"0840";
    tmp(08574) := x"0840";
    tmp(08575) := x"0020";
    tmp(08576) := x"0020";
    tmp(08577) := x"0020";
    tmp(08578) := x"0020";
    tmp(08579) := x"0020";
    tmp(08580) := x"0020";
    tmp(08581) := x"0020";
    tmp(08582) := x"0020";
    tmp(08583) := x"0020";
    tmp(08584) := x"0020";
    tmp(08585) := x"0020";
    tmp(08586) := x"0020";
    tmp(08587) := x"0020";
    tmp(08588) := x"0020";
    tmp(08589) := x"0020";
    tmp(08590) := x"0020";
    tmp(08591) := x"0020";
    tmp(08592) := x"0020";
    tmp(08593) := x"0020";
    tmp(08594) := x"0020";
    tmp(08595) := x"0020";
    tmp(08596) := x"0020";
    tmp(08597) := x"ffff";
    tmp(08598) := x"ffff";
    tmp(08599) := x"ffff";
    tmp(08600) := x"ffff";
    tmp(08601) := x"ffff";
    tmp(08602) := x"ffff";
    tmp(08603) := x"ffff";
    tmp(08604) := x"ffff";
    tmp(08605) := x"ffff";
    tmp(08606) := x"ffff";
    tmp(08607) := x"ffff";
    tmp(08608) := x"ffff";
    tmp(08609) := x"ffff";
    tmp(08610) := x"ffff";
    tmp(08611) := x"ffff";
    tmp(08612) := x"ffff";
    tmp(08613) := x"ffff";
    tmp(08614) := x"ffff";
    tmp(08615) := x"ffff";
    tmp(08616) := x"ffff";
    tmp(08617) := x"ffff";
    tmp(08618) := x"ffff";
    tmp(08619) := x"ffff";
    tmp(08620) := x"ffff";
    tmp(08621) := x"ffff";
    tmp(08622) := x"ffff";
    tmp(08623) := x"ffff";
    tmp(08624) := x"ffff";
    tmp(08625) := x"ffff";
    tmp(08626) := x"ffff";
    tmp(08627) := x"ffff";
    tmp(08628) := x"ffff";
    tmp(08629) := x"ffff";
    tmp(08630) := x"ffff";
    tmp(08631) := x"ffff";
    tmp(08632) := x"ffff";
    tmp(08633) := x"ffff";
    tmp(08634) := x"ffff";
    tmp(08635) := x"ffff";
    tmp(08636) := x"ffff";
    tmp(08637) := x"0820";
    tmp(08638) := x"0820";
    tmp(08639) := x"0820";
    tmp(08640) := x"0000";
    tmp(08641) := x"0040";
    tmp(08642) := x"0040";
    tmp(08643) := x"0040";
    tmp(08644) := x"0040";
    tmp(08645) := x"0040";
    tmp(08646) := x"0040";
    tmp(08647) := x"0040";
    tmp(08648) := x"0040";
    tmp(08649) := x"0040";
    tmp(08650) := x"0020";
    tmp(08651) := x"0020";
    tmp(08652) := x"0020";
    tmp(08653) := x"0020";
    tmp(08654) := x"0020";
    tmp(08655) := x"0020";
    tmp(08656) := x"0020";
    tmp(08657) := x"0020";
    tmp(08658) := x"0020";
    tmp(08659) := x"0020";
    tmp(08660) := x"0020";
    tmp(08661) := x"0020";
    tmp(08662) := x"0820";
    tmp(08663) := x"0820";
    tmp(08664) := x"0820";
    tmp(08665) := x"0820";
    tmp(08666) := x"0820";
    tmp(08667) := x"0820";
    tmp(08668) := x"0820";
    tmp(08669) := x"0820";
    tmp(08670) := x"0820";
    tmp(08671) := x"0820";
    tmp(08672) := x"0820";
    tmp(08673) := x"0820";
    tmp(08674) := x"0820";
    tmp(08675) := x"0820";
    tmp(08676) := x"0820";
    tmp(08677) := x"0820";
    tmp(08678) := x"0820";
    tmp(08679) := x"0820";
    tmp(08680) := x"0820";
    tmp(08681) := x"0820";
    tmp(08682) := x"0840";
    tmp(08683) := x"0840";
    tmp(08684) := x"0840";
    tmp(08685) := x"0840";
    tmp(08686) := x"0840";
    tmp(08687) := x"0840";
    tmp(08688) := x"0840";
    tmp(08689) := x"0840";
    tmp(08690) := x"0840";
    tmp(08691) := x"0840";
    tmp(08692) := x"0840";
    tmp(08693) := x"0840";
    tmp(08694) := x"0840";
    tmp(08695) := x"0840";
    tmp(08696) := x"0840";
    tmp(08697) := x"0840";
    tmp(08698) := x"0840";
    tmp(08699) := x"0840";
    tmp(08700) := x"0840";
    tmp(08701) := x"0840";
    tmp(08702) := x"0840";
    tmp(08703) := x"0840";
    tmp(08704) := x"0840";
    tmp(08705) := x"0840";
    tmp(08706) := x"0840";
    tmp(08707) := x"0841";
    tmp(08708) := x"0840";
    tmp(08709) := x"0841";
    tmp(08710) := x"0840";
    tmp(08711) := x"0840";
    tmp(08712) := x"0840";
    tmp(08713) := x"0840";
    tmp(08714) := x"0840";
    tmp(08715) := x"0840";
    tmp(08716) := x"0840";
    tmp(08717) := x"0840";
    tmp(08718) := x"0840";
    tmp(08719) := x"0840";
    tmp(08720) := x"0840";
    tmp(08721) := x"0840";
    tmp(08722) := x"0860";
    tmp(08723) := x"0860";
    tmp(08724) := x"0860";
    tmp(08725) := x"0860";
    tmp(08726) := x"0860";
    tmp(08727) := x"0860";
    tmp(08728) := x"0860";
    tmp(08729) := x"0860";
    tmp(08730) := x"0880";
    tmp(08731) := x"0880";
    tmp(08732) := x"0880";
    tmp(08733) := x"0880";
    tmp(08734) := x"0880";
    tmp(08735) := x"0880";
    tmp(08736) := x"0880";
    tmp(08737) := x"0880";
    tmp(08738) := x"0880";
    tmp(08739) := x"0880";
    tmp(08740) := x"0860";
    tmp(08741) := x"0000";
    tmp(08742) := x"0000";
    tmp(08743) := x"0000";
    tmp(08744) := x"0000";
    tmp(08745) := x"0000";
    tmp(08746) := x"0000";
    tmp(08747) := x"0000";
    tmp(08748) := x"0000";
    tmp(08749) := x"0000";
    tmp(08750) := x"0000";
    tmp(08751) := x"0000";
    tmp(08752) := x"0821";
    tmp(08753) := x"0020";
    tmp(08754) := x"0000";
    tmp(08755) := x"0000";
    tmp(08756) := x"0000";
    tmp(08757) := x"0000";
    tmp(08758) := x"0000";
    tmp(08759) := x"0020";
    tmp(08760) := x"0000";
    tmp(08761) := x"0000";
    tmp(08762) := x"0000";
    tmp(08763) := x"0000";
    tmp(08764) := x"0000";
    tmp(08765) := x"0000";
    tmp(08766) := x"0000";
    tmp(08767) := x"0000";
    tmp(08768) := x"0000";
    tmp(08769) := x"0020";
    tmp(08770) := x"0020";
    tmp(08771) := x"0000";
    tmp(08772) := x"0000";
    tmp(08773) := x"0020";
    tmp(08774) := x"0020";
    tmp(08775) := x"0000";
    tmp(08776) := x"0000";
    tmp(08777) := x"0020";
    tmp(08778) := x"0020";
    tmp(08779) := x"0821";
    tmp(08780) := x"0841";
    tmp(08781) := x"0821";
    tmp(08782) := x"0821";
    tmp(08783) := x"0821";
    tmp(08784) := x"0841";
    tmp(08785) := x"1061";
    tmp(08786) := x"18c2";
    tmp(08787) := x"18c2";
    tmp(08788) := x"10a1";
    tmp(08789) := x"08c0";
    tmp(08790) := x"08a0";
    tmp(08791) := x"08a0";
    tmp(08792) := x"08a0";
    tmp(08793) := x"08a0";
    tmp(08794) := x"08a0";
    tmp(08795) := x"08a0";
    tmp(08796) := x"08a0";
    tmp(08797) := x"08a0";
    tmp(08798) := x"08a0";
    tmp(08799) := x"0880";
    tmp(08800) := x"0880";
    tmp(08801) := x"0880";
    tmp(08802) := x"0880";
    tmp(08803) := x"0880";
    tmp(08804) := x"0880";
    tmp(08805) := x"0860";
    tmp(08806) := x"0860";
    tmp(08807) := x"0860";
    tmp(08808) := x"0860";
    tmp(08809) := x"0840";
    tmp(08810) := x"0840";
    tmp(08811) := x"0840";
    tmp(08812) := x"0840";
    tmp(08813) := x"0840";
    tmp(08814) := x"0840";
    tmp(08815) := x"0840";
    tmp(08816) := x"0020";
    tmp(08817) := x"0020";
    tmp(08818) := x"0020";
    tmp(08819) := x"0020";
    tmp(08820) := x"0020";
    tmp(08821) := x"0020";
    tmp(08822) := x"0020";
    tmp(08823) := x"0020";
    tmp(08824) := x"0020";
    tmp(08825) := x"0020";
    tmp(08826) := x"0020";
    tmp(08827) := x"0020";
    tmp(08828) := x"0020";
    tmp(08829) := x"0020";
    tmp(08830) := x"0020";
    tmp(08831) := x"0020";
    tmp(08832) := x"0020";
    tmp(08833) := x"0020";
    tmp(08834) := x"0020";
    tmp(08835) := x"0020";
    tmp(08836) := x"0020";
    tmp(08837) := x"ffff";
    tmp(08838) := x"ffff";
    tmp(08839) := x"ffff";
    tmp(08840) := x"ffff";
    tmp(08841) := x"ffff";
    tmp(08842) := x"ffff";
    tmp(08843) := x"ffff";
    tmp(08844) := x"ffff";
    tmp(08845) := x"ffff";
    tmp(08846) := x"ffff";
    tmp(08847) := x"ffff";
    tmp(08848) := x"ffff";
    tmp(08849) := x"ffff";
    tmp(08850) := x"ffff";
    tmp(08851) := x"ffff";
    tmp(08852) := x"ffff";
    tmp(08853) := x"ffff";
    tmp(08854) := x"ffff";
    tmp(08855) := x"ffff";
    tmp(08856) := x"ffff";
    tmp(08857) := x"ffff";
    tmp(08858) := x"ffff";
    tmp(08859) := x"ffff";
    tmp(08860) := x"ffff";
    tmp(08861) := x"ffff";
    tmp(08862) := x"ffff";
    tmp(08863) := x"ffff";
    tmp(08864) := x"ffff";
    tmp(08865) := x"ffff";
    tmp(08866) := x"ffff";
    tmp(08867) := x"ffff";
    tmp(08868) := x"ffff";
    tmp(08869) := x"ffff";
    tmp(08870) := x"ffff";
    tmp(08871) := x"ffff";
    tmp(08872) := x"ffff";
    tmp(08873) := x"ffff";
    tmp(08874) := x"ffff";
    tmp(08875) := x"ffff";
    tmp(08876) := x"ffff";
    tmp(08877) := x"0820";
    tmp(08878) := x"0820";
    tmp(08879) := x"0820";
    tmp(08880) := x"0000";
    tmp(08881) := x"0040";
    tmp(08882) := x"0040";
    tmp(08883) := x"0040";
    tmp(08884) := x"0040";
    tmp(08885) := x"0040";
    tmp(08886) := x"0040";
    tmp(08887) := x"0040";
    tmp(08888) := x"0040";
    tmp(08889) := x"0040";
    tmp(08890) := x"0020";
    tmp(08891) := x"0020";
    tmp(08892) := x"0020";
    tmp(08893) := x"0020";
    tmp(08894) := x"0020";
    tmp(08895) := x"0020";
    tmp(08896) := x"0020";
    tmp(08897) := x"0020";
    tmp(08898) := x"0020";
    tmp(08899) := x"0020";
    tmp(08900) := x"0020";
    tmp(08901) := x"0020";
    tmp(08902) := x"0020";
    tmp(08903) := x"0820";
    tmp(08904) := x"0820";
    tmp(08905) := x"0820";
    tmp(08906) := x"0820";
    tmp(08907) := x"0820";
    tmp(08908) := x"0820";
    tmp(08909) := x"0820";
    tmp(08910) := x"0820";
    tmp(08911) := x"0820";
    tmp(08912) := x"0820";
    tmp(08913) := x"0820";
    tmp(08914) := x"0820";
    tmp(08915) := x"0820";
    tmp(08916) := x"0820";
    tmp(08917) := x"0820";
    tmp(08918) := x"0820";
    tmp(08919) := x"0820";
    tmp(08920) := x"0820";
    tmp(08921) := x"0820";
    tmp(08922) := x"0820";
    tmp(08923) := x"0840";
    tmp(08924) := x"0820";
    tmp(08925) := x"0840";
    tmp(08926) := x"0840";
    tmp(08927) := x"0840";
    tmp(08928) := x"0840";
    tmp(08929) := x"0840";
    tmp(08930) := x"0840";
    tmp(08931) := x"0840";
    tmp(08932) := x"0840";
    tmp(08933) := x"0840";
    tmp(08934) := x"0840";
    tmp(08935) := x"0840";
    tmp(08936) := x"0840";
    tmp(08937) := x"0840";
    tmp(08938) := x"0840";
    tmp(08939) := x"0840";
    tmp(08940) := x"0840";
    tmp(08941) := x"0840";
    tmp(08942) := x"0840";
    tmp(08943) := x"0840";
    tmp(08944) := x"0840";
    tmp(08945) := x"0840";
    tmp(08946) := x"0840";
    tmp(08947) := x"0840";
    tmp(08948) := x"0840";
    tmp(08949) := x"0840";
    tmp(08950) := x"0840";
    tmp(08951) := x"0840";
    tmp(08952) := x"0841";
    tmp(08953) := x"0841";
    tmp(08954) := x"0840";
    tmp(08955) := x"0840";
    tmp(08956) := x"0840";
    tmp(08957) := x"0840";
    tmp(08958) := x"0840";
    tmp(08959) := x"0840";
    tmp(08960) := x"0840";
    tmp(08961) := x"0860";
    tmp(08962) := x"0860";
    tmp(08963) := x"0860";
    tmp(08964) := x"0860";
    tmp(08965) := x"0860";
    tmp(08966) := x"0860";
    tmp(08967) := x"0860";
    tmp(08968) := x"0860";
    tmp(08969) := x"0860";
    tmp(08970) := x"0880";
    tmp(08971) := x"0880";
    tmp(08972) := x"0880";
    tmp(08973) := x"0880";
    tmp(08974) := x"0880";
    tmp(08975) := x"0880";
    tmp(08976) := x"0880";
    tmp(08977) := x"0880";
    tmp(08978) := x"0860";
    tmp(08979) := x"0880";
    tmp(08980) := x"0840";
    tmp(08981) := x"0000";
    tmp(08982) := x"0000";
    tmp(08983) := x"0000";
    tmp(08984) := x"0000";
    tmp(08985) := x"0000";
    tmp(08986) := x"0000";
    tmp(08987) := x"0000";
    tmp(08988) := x"0000";
    tmp(08989) := x"0000";
    tmp(08990) := x"0000";
    tmp(08991) := x"0000";
    tmp(08992) := x"0821";
    tmp(08993) := x"0821";
    tmp(08994) := x"0000";
    tmp(08995) := x"0000";
    tmp(08996) := x"0000";
    tmp(08997) := x"0000";
    tmp(08998) := x"0000";
    tmp(08999) := x"0000";
    tmp(09000) := x"0000";
    tmp(09001) := x"0000";
    tmp(09002) := x"0000";
    tmp(09003) := x"0000";
    tmp(09004) := x"0000";
    tmp(09005) := x"0000";
    tmp(09006) := x"0000";
    tmp(09007) := x"0000";
    tmp(09008) := x"0000";
    tmp(09009) := x"0020";
    tmp(09010) := x"0020";
    tmp(09011) := x"0020";
    tmp(09012) := x"0000";
    tmp(09013) := x"0000";
    tmp(09014) := x"0020";
    tmp(09015) := x"0020";
    tmp(09016) := x"0821";
    tmp(09017) := x"0821";
    tmp(09018) := x"0821";
    tmp(09019) := x"0841";
    tmp(09020) := x"0841";
    tmp(09021) := x"0841";
    tmp(09022) := x"0841";
    tmp(09023) := x"0821";
    tmp(09024) := x"0841";
    tmp(09025) := x"0841";
    tmp(09026) := x"18a2";
    tmp(09027) := x"20e2";
    tmp(09028) := x"1081";
    tmp(09029) := x"10c1";
    tmp(09030) := x"08a0";
    tmp(09031) := x"08a0";
    tmp(09032) := x"08c0";
    tmp(09033) := x"08c0";
    tmp(09034) := x"08c0";
    tmp(09035) := x"08c0";
    tmp(09036) := x"08c0";
    tmp(09037) := x"08a0";
    tmp(09038) := x"08a0";
    tmp(09039) := x"08a0";
    tmp(09040) := x"08a0";
    tmp(09041) := x"08a0";
    tmp(09042) := x"08a0";
    tmp(09043) := x"0880";
    tmp(09044) := x"0880";
    tmp(09045) := x"0880";
    tmp(09046) := x"0880";
    tmp(09047) := x"0880";
    tmp(09048) := x"0860";
    tmp(09049) := x"0860";
    tmp(09050) := x"0860";
    tmp(09051) := x"0860";
    tmp(09052) := x"0840";
    tmp(09053) := x"0840";
    tmp(09054) := x"0840";
    tmp(09055) := x"0840";
    tmp(09056) := x"0840";
    tmp(09057) := x"0840";
    tmp(09058) := x"0020";
    tmp(09059) := x"0020";
    tmp(09060) := x"0020";
    tmp(09061) := x"0020";
    tmp(09062) := x"0020";
    tmp(09063) := x"0020";
    tmp(09064) := x"0020";
    tmp(09065) := x"0020";
    tmp(09066) := x"0020";
    tmp(09067) := x"0020";
    tmp(09068) := x"0020";
    tmp(09069) := x"0020";
    tmp(09070) := x"0020";
    tmp(09071) := x"0020";
    tmp(09072) := x"0020";
    tmp(09073) := x"0020";
    tmp(09074) := x"0020";
    tmp(09075) := x"0000";
    tmp(09076) := x"0020";
    tmp(09077) := x"ffff";
    tmp(09078) := x"ffff";
    tmp(09079) := x"ffff";
    tmp(09080) := x"ffff";
    tmp(09081) := x"ffff";
    tmp(09082) := x"ffff";
    tmp(09083) := x"ffff";
    tmp(09084) := x"ffff";
    tmp(09085) := x"ffff";
    tmp(09086) := x"ffff";
    tmp(09087) := x"ffff";
    tmp(09088) := x"ffff";
    tmp(09089) := x"ffff";
    tmp(09090) := x"ffff";
    tmp(09091) := x"ffff";
    tmp(09092) := x"ffff";
    tmp(09093) := x"ffff";
    tmp(09094) := x"ffff";
    tmp(09095) := x"ffff";
    tmp(09096) := x"ffff";
    tmp(09097) := x"ffff";
    tmp(09098) := x"ffff";
    tmp(09099) := x"ffff";
    tmp(09100) := x"ffff";
    tmp(09101) := x"ffff";
    tmp(09102) := x"ffff";
    tmp(09103) := x"ffff";
    tmp(09104) := x"ffff";
    tmp(09105) := x"ffff";
    tmp(09106) := x"ffff";
    tmp(09107) := x"ffff";
    tmp(09108) := x"ffff";
    tmp(09109) := x"ffff";
    tmp(09110) := x"ffff";
    tmp(09111) := x"ffff";
    tmp(09112) := x"ffff";
    tmp(09113) := x"ffff";
    tmp(09114) := x"ffff";
    tmp(09115) := x"ffff";
    tmp(09116) := x"ffff";
    tmp(09117) := x"0820";
    tmp(09118) := x"0820";
    tmp(09119) := x"0820";
    tmp(09120) := x"0000";
    tmp(09121) := x"0040";
    tmp(09122) := x"0040";
    tmp(09123) := x"0040";
    tmp(09124) := x"0040";
    tmp(09125) := x"0040";
    tmp(09126) := x"0040";
    tmp(09127) := x"0040";
    tmp(09128) := x"0040";
    tmp(09129) := x"0020";
    tmp(09130) := x"0020";
    tmp(09131) := x"0020";
    tmp(09132) := x"0020";
    tmp(09133) := x"0020";
    tmp(09134) := x"0020";
    tmp(09135) := x"0020";
    tmp(09136) := x"0020";
    tmp(09137) := x"0020";
    tmp(09138) := x"0020";
    tmp(09139) := x"0020";
    tmp(09140) := x"0020";
    tmp(09141) := x"0020";
    tmp(09142) := x"0820";
    tmp(09143) := x"0820";
    tmp(09144) := x"0820";
    tmp(09145) := x"0820";
    tmp(09146) := x"0820";
    tmp(09147) := x"0820";
    tmp(09148) := x"0820";
    tmp(09149) := x"0820";
    tmp(09150) := x"0820";
    tmp(09151) := x"0820";
    tmp(09152) := x"0820";
    tmp(09153) := x"0820";
    tmp(09154) := x"0820";
    tmp(09155) := x"0820";
    tmp(09156) := x"0820";
    tmp(09157) := x"0820";
    tmp(09158) := x"0820";
    tmp(09159) := x"0820";
    tmp(09160) := x"0820";
    tmp(09161) := x"0820";
    tmp(09162) := x"0820";
    tmp(09163) := x"0820";
    tmp(09164) := x"0840";
    tmp(09165) := x"0840";
    tmp(09166) := x"0820";
    tmp(09167) := x"0840";
    tmp(09168) := x"0840";
    tmp(09169) := x"0840";
    tmp(09170) := x"0840";
    tmp(09171) := x"0840";
    tmp(09172) := x"0840";
    tmp(09173) := x"0840";
    tmp(09174) := x"0840";
    tmp(09175) := x"0840";
    tmp(09176) := x"0840";
    tmp(09177) := x"0840";
    tmp(09178) := x"0840";
    tmp(09179) := x"0840";
    tmp(09180) := x"0840";
    tmp(09181) := x"0840";
    tmp(09182) := x"0840";
    tmp(09183) := x"0840";
    tmp(09184) := x"0840";
    tmp(09185) := x"0840";
    tmp(09186) := x"0840";
    tmp(09187) := x"0840";
    tmp(09188) := x"0841";
    tmp(09189) := x"0840";
    tmp(09190) := x"0840";
    tmp(09191) := x"0841";
    tmp(09192) := x"0840";
    tmp(09193) := x"0840";
    tmp(09194) := x"0840";
    tmp(09195) := x"0840";
    tmp(09196) := x"0840";
    tmp(09197) := x"0840";
    tmp(09198) := x"0840";
    tmp(09199) := x"0840";
    tmp(09200) := x"0840";
    tmp(09201) := x"0860";
    tmp(09202) := x"0860";
    tmp(09203) := x"0860";
    tmp(09204) := x"0860";
    tmp(09205) := x"0860";
    tmp(09206) := x"0860";
    tmp(09207) := x"0860";
    tmp(09208) := x"0860";
    tmp(09209) := x"0860";
    tmp(09210) := x"0880";
    tmp(09211) := x"0880";
    tmp(09212) := x"0880";
    tmp(09213) := x"0880";
    tmp(09214) := x"0880";
    tmp(09215) := x"0880";
    tmp(09216) := x"0880";
    tmp(09217) := x"0860";
    tmp(09218) := x"0860";
    tmp(09219) := x"0880";
    tmp(09220) := x"0020";
    tmp(09221) := x"0000";
    tmp(09222) := x"0000";
    tmp(09223) := x"0000";
    tmp(09224) := x"0000";
    tmp(09225) := x"0000";
    tmp(09226) := x"0000";
    tmp(09227) := x"0000";
    tmp(09228) := x"0000";
    tmp(09229) := x"0000";
    tmp(09230) := x"0000";
    tmp(09231) := x"0000";
    tmp(09232) := x"0000";
    tmp(09233) := x"0841";
    tmp(09234) := x"0000";
    tmp(09235) := x"0000";
    tmp(09236) := x"0000";
    tmp(09237) := x"0000";
    tmp(09238) := x"0020";
    tmp(09239) := x"0000";
    tmp(09240) := x"0000";
    tmp(09241) := x"0000";
    tmp(09242) := x"0000";
    tmp(09243) := x"0000";
    tmp(09244) := x"0000";
    tmp(09245) := x"0000";
    tmp(09246) := x"0000";
    tmp(09247) := x"0000";
    tmp(09248) := x"0000";
    tmp(09249) := x"0000";
    tmp(09250) := x"0000";
    tmp(09251) := x"0020";
    tmp(09252) := x"0020";
    tmp(09253) := x"0020";
    tmp(09254) := x"0020";
    tmp(09255) := x"0020";
    tmp(09256) := x"0020";
    tmp(09257) := x"0020";
    tmp(09258) := x"0821";
    tmp(09259) := x"0021";
    tmp(09260) := x"0841";
    tmp(09261) := x"0841";
    tmp(09262) := x"0821";
    tmp(09263) := x"0020";
    tmp(09264) := x"0821";
    tmp(09265) := x"0841";
    tmp(09266) := x"1081";
    tmp(09267) := x"2102";
    tmp(09268) := x"20e2";
    tmp(09269) := x"10a1";
    tmp(09270) := x"10c0";
    tmp(09271) := x"08a0";
    tmp(09272) := x"08c0";
    tmp(09273) := x"08c0";
    tmp(09274) := x"08c0";
    tmp(09275) := x"08c0";
    tmp(09276) := x"08c0";
    tmp(09277) := x"08c0";
    tmp(09278) := x"08c0";
    tmp(09279) := x"08c0";
    tmp(09280) := x"08c0";
    tmp(09281) := x"08a0";
    tmp(09282) := x"08a0";
    tmp(09283) := x"08a0";
    tmp(09284) := x"08a0";
    tmp(09285) := x"0880";
    tmp(09286) := x"0880";
    tmp(09287) := x"0880";
    tmp(09288) := x"0880";
    tmp(09289) := x"0880";
    tmp(09290) := x"0880";
    tmp(09291) := x"0860";
    tmp(09292) := x"0860";
    tmp(09293) := x"0860";
    tmp(09294) := x"0860";
    tmp(09295) := x"0860";
    tmp(09296) := x"0840";
    tmp(09297) := x"0840";
    tmp(09298) := x"0840";
    tmp(09299) := x"0040";
    tmp(09300) := x"0040";
    tmp(09301) := x"0020";
    tmp(09302) := x"0020";
    tmp(09303) := x"0020";
    tmp(09304) := x"0020";
    tmp(09305) := x"0020";
    tmp(09306) := x"0020";
    tmp(09307) := x"0020";
    tmp(09308) := x"0020";
    tmp(09309) := x"0020";
    tmp(09310) := x"0000";
    tmp(09311) := x"0000";
    tmp(09312) := x"0000";
    tmp(09313) := x"0000";
    tmp(09314) := x"0000";
    tmp(09315) := x"0000";
    tmp(09316) := x"0000";
    tmp(09317) := x"ffff";
    tmp(09318) := x"ffff";
    tmp(09319) := x"ffff";
    tmp(09320) := x"ffff";
    tmp(09321) := x"ffff";
    tmp(09322) := x"ffff";
    tmp(09323) := x"ffff";
    tmp(09324) := x"ffff";
    tmp(09325) := x"ffff";
    tmp(09326) := x"ffff";
    tmp(09327) := x"ffff";
    tmp(09328) := x"ffff";
    tmp(09329) := x"ffff";
    tmp(09330) := x"ffff";
    tmp(09331) := x"ffff";
    tmp(09332) := x"ffff";
    tmp(09333) := x"ffff";
    tmp(09334) := x"ffff";
    tmp(09335) := x"ffff";
    tmp(09336) := x"ffff";
    tmp(09337) := x"ffff";
    tmp(09338) := x"ffff";
    tmp(09339) := x"ffff";
    tmp(09340) := x"ffff";
    tmp(09341) := x"ffff";
    tmp(09342) := x"ffff";
    tmp(09343) := x"ffff";
    tmp(09344) := x"ffff";
    tmp(09345) := x"ffff";
    tmp(09346) := x"ffff";
    tmp(09347) := x"ffff";
    tmp(09348) := x"ffff";
    tmp(09349) := x"ffff";
    tmp(09350) := x"ffff";
    tmp(09351) := x"ffff";
    tmp(09352) := x"ffff";
    tmp(09353) := x"ffff";
    tmp(09354) := x"ffff";
    tmp(09355) := x"ffff";
    tmp(09356) := x"ffff";
    tmp(09357) := x"0820";
    tmp(09358) := x"0820";
    tmp(09359) := x"0820";
    tmp(09360) := x"0000";
    tmp(09361) := x"0040";
    tmp(09362) := x"0040";
    tmp(09363) := x"0040";
    tmp(09364) := x"0040";
    tmp(09365) := x"0040";
    tmp(09366) := x"0040";
    tmp(09367) := x"0040";
    tmp(09368) := x"0020";
    tmp(09369) := x"0020";
    tmp(09370) := x"0020";
    tmp(09371) := x"0020";
    tmp(09372) := x"0020";
    tmp(09373) := x"0020";
    tmp(09374) := x"0020";
    tmp(09375) := x"0020";
    tmp(09376) := x"0020";
    tmp(09377) := x"0020";
    tmp(09378) := x"0020";
    tmp(09379) := x"0020";
    tmp(09380) := x"0020";
    tmp(09381) := x"0820";
    tmp(09382) := x"0820";
    tmp(09383) := x"0820";
    tmp(09384) := x"0820";
    tmp(09385) := x"0820";
    tmp(09386) := x"0820";
    tmp(09387) := x"0820";
    tmp(09388) := x"0820";
    tmp(09389) := x"0820";
    tmp(09390) := x"0820";
    tmp(09391) := x"0820";
    tmp(09392) := x"0820";
    tmp(09393) := x"0820";
    tmp(09394) := x"0820";
    tmp(09395) := x"0820";
    tmp(09396) := x"0820";
    tmp(09397) := x"0820";
    tmp(09398) := x"0820";
    tmp(09399) := x"0820";
    tmp(09400) := x"0820";
    tmp(09401) := x"0820";
    tmp(09402) := x"0820";
    tmp(09403) := x"0840";
    tmp(09404) := x"0840";
    tmp(09405) := x"0840";
    tmp(09406) := x"0840";
    tmp(09407) := x"0840";
    tmp(09408) := x"0840";
    tmp(09409) := x"0840";
    tmp(09410) := x"0840";
    tmp(09411) := x"0840";
    tmp(09412) := x"0840";
    tmp(09413) := x"0840";
    tmp(09414) := x"0840";
    tmp(09415) := x"0840";
    tmp(09416) := x"0840";
    tmp(09417) := x"0840";
    tmp(09418) := x"0840";
    tmp(09419) := x"0840";
    tmp(09420) := x"0840";
    tmp(09421) := x"0840";
    tmp(09422) := x"0840";
    tmp(09423) := x"0840";
    tmp(09424) := x"0840";
    tmp(09425) := x"0840";
    tmp(09426) := x"0840";
    tmp(09427) := x"0840";
    tmp(09428) := x"0841";
    tmp(09429) := x"0840";
    tmp(09430) := x"0840";
    tmp(09431) := x"0840";
    tmp(09432) := x"0840";
    tmp(09433) := x"0840";
    tmp(09434) := x"0840";
    tmp(09435) := x"0840";
    tmp(09436) := x"0840";
    tmp(09437) := x"0840";
    tmp(09438) := x"0840";
    tmp(09439) := x"0840";
    tmp(09440) := x"0840";
    tmp(09441) := x"0840";
    tmp(09442) := x"0840";
    tmp(09443) := x"0860";
    tmp(09444) := x"0860";
    tmp(09445) := x"0860";
    tmp(09446) := x"0860";
    tmp(09447) := x"0860";
    tmp(09448) := x"0860";
    tmp(09449) := x"0880";
    tmp(09450) := x"0880";
    tmp(09451) := x"0880";
    tmp(09452) := x"0880";
    tmp(09453) := x"0880";
    tmp(09454) := x"0880";
    tmp(09455) := x"0880";
    tmp(09456) := x"0880";
    tmp(09457) := x"0860";
    tmp(09458) := x"0860";
    tmp(09459) := x"0860";
    tmp(09460) := x"0020";
    tmp(09461) := x"0000";
    tmp(09462) := x"0000";
    tmp(09463) := x"0000";
    tmp(09464) := x"0000";
    tmp(09465) := x"0000";
    tmp(09466) := x"0000";
    tmp(09467) := x"0000";
    tmp(09468) := x"0000";
    tmp(09469) := x"0000";
    tmp(09470) := x"0000";
    tmp(09471) := x"0000";
    tmp(09472) := x"0000";
    tmp(09473) := x"0000";
    tmp(09474) := x"0020";
    tmp(09475) := x"0000";
    tmp(09476) := x"0000";
    tmp(09477) := x"0000";
    tmp(09478) := x"0020";
    tmp(09479) := x"0000";
    tmp(09480) := x"0000";
    tmp(09481) := x"0000";
    tmp(09482) := x"0000";
    tmp(09483) := x"0000";
    tmp(09484) := x"0000";
    tmp(09485) := x"0000";
    tmp(09486) := x"0000";
    tmp(09487) := x"0000";
    tmp(09488) := x"0000";
    tmp(09489) := x"0000";
    tmp(09490) := x"0000";
    tmp(09491) := x"0000";
    tmp(09492) := x"0821";
    tmp(09493) := x"0020";
    tmp(09494) := x"0000";
    tmp(09495) := x"0020";
    tmp(09496) := x"0020";
    tmp(09497) := x"0020";
    tmp(09498) := x"0821";
    tmp(09499) := x"0020";
    tmp(09500) := x"0821";
    tmp(09501) := x"0841";
    tmp(09502) := x"0841";
    tmp(09503) := x"0821";
    tmp(09504) := x"0821";
    tmp(09505) := x"0821";
    tmp(09506) := x"0861";
    tmp(09507) := x"20e2";
    tmp(09508) := x"3143";
    tmp(09509) := x"10a1";
    tmp(09510) := x"31a3";
    tmp(09511) := x"1921";
    tmp(09512) := x"10c0";
    tmp(09513) := x"08c0";
    tmp(09514) := x"08c0";
    tmp(09515) := x"08e0";
    tmp(09516) := x"08c0";
    tmp(09517) := x"08c0";
    tmp(09518) := x"08e0";
    tmp(09519) := x"08e0";
    tmp(09520) := x"08c0";
    tmp(09521) := x"08c0";
    tmp(09522) := x"08c0";
    tmp(09523) := x"08c0";
    tmp(09524) := x"08a0";
    tmp(09525) := x"08a0";
    tmp(09526) := x"08a0";
    tmp(09527) := x"08a0";
    tmp(09528) := x"08a0";
    tmp(09529) := x"08a0";
    tmp(09530) := x"0880";
    tmp(09531) := x"0880";
    tmp(09532) := x"0880";
    tmp(09533) := x"0880";
    tmp(09534) := x"0860";
    tmp(09535) := x"0860";
    tmp(09536) := x"0860";
    tmp(09537) := x"0860";
    tmp(09538) := x"0860";
    tmp(09539) := x"0840";
    tmp(09540) := x"0040";
    tmp(09541) := x"0040";
    tmp(09542) := x"0040";
    tmp(09543) := x"0040";
    tmp(09544) := x"0020";
    tmp(09545) := x"0020";
    tmp(09546) := x"0020";
    tmp(09547) := x"0020";
    tmp(09548) := x"0020";
    tmp(09549) := x"0020";
    tmp(09550) := x"0020";
    tmp(09551) := x"0020";
    tmp(09552) := x"0000";
    tmp(09553) := x"0000";
    tmp(09554) := x"0000";
    tmp(09555) := x"0000";
    tmp(09556) := x"0000";
    tmp(09557) := x"ffff";
    tmp(09558) := x"ffff";
    tmp(09559) := x"ffff";
    tmp(09560) := x"ffff";
    tmp(09561) := x"ffff";
    tmp(09562) := x"ffff";
    tmp(09563) := x"ffff";
    tmp(09564) := x"ffff";
    tmp(09565) := x"ffff";
    tmp(09566) := x"ffff";
    tmp(09567) := x"ffff";
    tmp(09568) := x"ffff";
    tmp(09569) := x"ffff";
    tmp(09570) := x"ffff";
    tmp(09571) := x"ffff";
    tmp(09572) := x"ffff";
    tmp(09573) := x"ffff";
    tmp(09574) := x"ffff";
    tmp(09575) := x"ffff";
    tmp(09576) := x"ffff";
    tmp(09577) := x"ffff";
    tmp(09578) := x"ffff";
    tmp(09579) := x"ffff";
    tmp(09580) := x"ffff";
    tmp(09581) := x"ffff";
    tmp(09582) := x"ffff";
    tmp(09583) := x"ffff";
    tmp(09584) := x"ffff";
    tmp(09585) := x"ffff";
    tmp(09586) := x"ffff";
    tmp(09587) := x"ffff";
    tmp(09588) := x"ffff";
    tmp(09589) := x"ffff";
    tmp(09590) := x"ffff";
    tmp(09591) := x"ffff";
    tmp(09592) := x"ffff";
    tmp(09593) := x"ffff";
    tmp(09594) := x"ffff";
    tmp(09595) := x"ffff";
    tmp(09596) := x"ffff";
    tmp(09597) := x"0820";
    tmp(09598) := x"0820";
    tmp(09599) := x"0820";
    tmp(09600) := x"0000";
    tmp(09601) := x"08a1";
    tmp(09602) := x"0881";
    tmp(09603) := x"0881";
    tmp(09604) := x"0861";
    tmp(09605) := x"0861";
    tmp(09606) := x"0060";
    tmp(09607) := x"0040";
    tmp(09608) := x"0040";
    tmp(09609) := x"0020";
    tmp(09610) := x"0020";
    tmp(09611) := x"0020";
    tmp(09612) := x"0020";
    tmp(09613) := x"0020";
    tmp(09614) := x"0020";
    tmp(09615) := x"0020";
    tmp(09616) := x"0020";
    tmp(09617) := x"0020";
    tmp(09618) := x"0020";
    tmp(09619) := x"0020";
    tmp(09620) := x"0020";
    tmp(09621) := x"0020";
    tmp(09622) := x"0020";
    tmp(09623) := x"0820";
    tmp(09624) := x"0820";
    tmp(09625) := x"0820";
    tmp(09626) := x"0820";
    tmp(09627) := x"0820";
    tmp(09628) := x"0820";
    tmp(09629) := x"0820";
    tmp(09630) := x"0820";
    tmp(09631) := x"0820";
    tmp(09632) := x"0820";
    tmp(09633) := x"0820";
    tmp(09634) := x"0820";
    tmp(09635) := x"0820";
    tmp(09636) := x"0820";
    tmp(09637) := x"0820";
    tmp(09638) := x"0820";
    tmp(09639) := x"0820";
    tmp(09640) := x"0820";
    tmp(09641) := x"0820";
    tmp(09642) := x"0820";
    tmp(09643) := x"0820";
    tmp(09644) := x"0840";
    tmp(09645) := x"0820";
    tmp(09646) := x"0840";
    tmp(09647) := x"0840";
    tmp(09648) := x"0840";
    tmp(09649) := x"0820";
    tmp(09650) := x"0840";
    tmp(09651) := x"0840";
    tmp(09652) := x"0840";
    tmp(09653) := x"0840";
    tmp(09654) := x"0840";
    tmp(09655) := x"0840";
    tmp(09656) := x"0840";
    tmp(09657) := x"0840";
    tmp(09658) := x"0840";
    tmp(09659) := x"0840";
    tmp(09660) := x"0840";
    tmp(09661) := x"0840";
    tmp(09662) := x"0840";
    tmp(09663) := x"0840";
    tmp(09664) := x"0840";
    tmp(09665) := x"0840";
    tmp(09666) := x"0840";
    tmp(09667) := x"0840";
    tmp(09668) := x"0840";
    tmp(09669) := x"0840";
    tmp(09670) := x"0840";
    tmp(09671) := x"0840";
    tmp(09672) := x"0840";
    tmp(09673) := x"0840";
    tmp(09674) := x"0840";
    tmp(09675) := x"0840";
    tmp(09676) := x"0840";
    tmp(09677) := x"0840";
    tmp(09678) := x"0840";
    tmp(09679) := x"0840";
    tmp(09680) := x"0840";
    tmp(09681) := x"0840";
    tmp(09682) := x"0840";
    tmp(09683) := x"0840";
    tmp(09684) := x"0860";
    tmp(09685) := x"0860";
    tmp(09686) := x"0860";
    tmp(09687) := x"0860";
    tmp(09688) := x"0860";
    tmp(09689) := x"0880";
    tmp(09690) := x"0880";
    tmp(09691) := x"0880";
    tmp(09692) := x"0880";
    tmp(09693) := x"0880";
    tmp(09694) := x"0880";
    tmp(09695) := x"0880";
    tmp(09696) := x"0880";
    tmp(09697) := x"0860";
    tmp(09698) := x"0860";
    tmp(09699) := x"0840";
    tmp(09700) := x"0000";
    tmp(09701) := x"0000";
    tmp(09702) := x"0000";
    tmp(09703) := x"0000";
    tmp(09704) := x"0000";
    tmp(09705) := x"0000";
    tmp(09706) := x"0000";
    tmp(09707) := x"0000";
    tmp(09708) := x"0000";
    tmp(09709) := x"0000";
    tmp(09710) := x"0000";
    tmp(09711) := x"0000";
    tmp(09712) := x"0000";
    tmp(09713) := x"0000";
    tmp(09714) := x"0000";
    tmp(09715) := x"0841";
    tmp(09716) := x"0020";
    tmp(09717) := x"0000";
    tmp(09718) := x"0020";
    tmp(09719) := x"0000";
    tmp(09720) := x"0000";
    tmp(09721) := x"0000";
    tmp(09722) := x"0000";
    tmp(09723) := x"0000";
    tmp(09724) := x"0000";
    tmp(09725) := x"0020";
    tmp(09726) := x"0000";
    tmp(09727) := x"0000";
    tmp(09728) := x"0000";
    tmp(09729) := x"0000";
    tmp(09730) := x"0000";
    tmp(09731) := x"0000";
    tmp(09732) := x"0020";
    tmp(09733) := x"0020";
    tmp(09734) := x"0020";
    tmp(09735) := x"0000";
    tmp(09736) := x"0021";
    tmp(09737) := x"0020";
    tmp(09738) := x"0020";
    tmp(09739) := x"0020";
    tmp(09740) := x"0020";
    tmp(09741) := x"0821";
    tmp(09742) := x"0841";
    tmp(09743) := x"0821";
    tmp(09744) := x"0020";
    tmp(09745) := x"0820";
    tmp(09746) := x"0841";
    tmp(09747) := x"18c2";
    tmp(09748) := x"3143";
    tmp(09749) := x"20c2";
    tmp(09750) := x"49c5";
    tmp(09751) := x"d694";
    tmp(09752) := x"18e1";
    tmp(09753) := x"0880";
    tmp(09754) := x"08c0";
    tmp(09755) := x"08c0";
    tmp(09756) := x"08c0";
    tmp(09757) := x"08c0";
    tmp(09758) := x"08c0";
    tmp(09759) := x"08c0";
    tmp(09760) := x"08e0";
    tmp(09761) := x"08c0";
    tmp(09762) := x"08c0";
    tmp(09763) := x"08c0";
    tmp(09764) := x"08c0";
    tmp(09765) := x"08c0";
    tmp(09766) := x"08c0";
    tmp(09767) := x"08c0";
    tmp(09768) := x"08a0";
    tmp(09769) := x"08a0";
    tmp(09770) := x"08a0";
    tmp(09771) := x"08a0";
    tmp(09772) := x"08a0";
    tmp(09773) := x"0880";
    tmp(09774) := x"0880";
    tmp(09775) := x"0880";
    tmp(09776) := x"0860";
    tmp(09777) := x"0860";
    tmp(09778) := x"0860";
    tmp(09779) := x"0860";
    tmp(09780) := x"0860";
    tmp(09781) := x"0040";
    tmp(09782) := x"0040";
    tmp(09783) := x"0040";
    tmp(09784) := x"0040";
    tmp(09785) := x"0040";
    tmp(09786) := x"0020";
    tmp(09787) := x"0020";
    tmp(09788) := x"0020";
    tmp(09789) := x"0020";
    tmp(09790) := x"0020";
    tmp(09791) := x"0020";
    tmp(09792) := x"0020";
    tmp(09793) := x"0000";
    tmp(09794) := x"0000";
    tmp(09795) := x"0000";
    tmp(09796) := x"0000";
    tmp(09797) := x"ffff";
    tmp(09798) := x"ffff";
    tmp(09799) := x"ffff";
    tmp(09800) := x"ffff";
    tmp(09801) := x"ffff";
    tmp(09802) := x"ffff";
    tmp(09803) := x"ffff";
    tmp(09804) := x"ffff";
    tmp(09805) := x"ffff";
    tmp(09806) := x"ffff";
    tmp(09807) := x"ffff";
    tmp(09808) := x"ffff";
    tmp(09809) := x"ffff";
    tmp(09810) := x"ffff";
    tmp(09811) := x"ffff";
    tmp(09812) := x"ffff";
    tmp(09813) := x"ffff";
    tmp(09814) := x"ffff";
    tmp(09815) := x"ffff";
    tmp(09816) := x"ffff";
    tmp(09817) := x"ffff";
    tmp(09818) := x"ffff";
    tmp(09819) := x"ffff";
    tmp(09820) := x"ffff";
    tmp(09821) := x"ffff";
    tmp(09822) := x"ffff";
    tmp(09823) := x"ffff";
    tmp(09824) := x"ffff";
    tmp(09825) := x"ffff";
    tmp(09826) := x"ffff";
    tmp(09827) := x"ffff";
    tmp(09828) := x"ffff";
    tmp(09829) := x"ffff";
    tmp(09830) := x"ffff";
    tmp(09831) := x"ffff";
    tmp(09832) := x"ffff";
    tmp(09833) := x"ffff";
    tmp(09834) := x"ffff";
    tmp(09835) := x"ffff";
    tmp(09836) := x"ffff";
    tmp(09837) := x"0820";
    tmp(09838) := x"0820";
    tmp(09839) := x"0820";
    tmp(09840) := x"0000";
    tmp(09841) := x"0020";
    tmp(09842) := x"0020";
    tmp(09843) := x"0041";
    tmp(09844) := x"0041";
    tmp(09845) := x"0041";
    tmp(09846) := x"0862";
    tmp(09847) := x"0882";
    tmp(09848) := x"0882";
    tmp(09849) := x"0861";
    tmp(09850) := x"0861";
    tmp(09851) := x"0861";
    tmp(09852) := x"0861";
    tmp(09853) := x"0841";
    tmp(09854) := x"0040";
    tmp(09855) := x"0020";
    tmp(09856) := x"0020";
    tmp(09857) := x"0020";
    tmp(09858) := x"0020";
    tmp(09859) := x"0020";
    tmp(09860) := x"0020";
    tmp(09861) := x"0020";
    tmp(09862) := x"0020";
    tmp(09863) := x"0820";
    tmp(09864) := x"0820";
    tmp(09865) := x"0820";
    tmp(09866) := x"0820";
    tmp(09867) := x"0820";
    tmp(09868) := x"0820";
    tmp(09869) := x"0820";
    tmp(09870) := x"0820";
    tmp(09871) := x"0820";
    tmp(09872) := x"0820";
    tmp(09873) := x"0820";
    tmp(09874) := x"0820";
    tmp(09875) := x"0820";
    tmp(09876) := x"0820";
    tmp(09877) := x"0820";
    tmp(09878) := x"0820";
    tmp(09879) := x"0820";
    tmp(09880) := x"0820";
    tmp(09881) := x"0820";
    tmp(09882) := x"0820";
    tmp(09883) := x"0840";
    tmp(09884) := x"0820";
    tmp(09885) := x"0820";
    tmp(09886) := x"0840";
    tmp(09887) := x"0820";
    tmp(09888) := x"0820";
    tmp(09889) := x"0840";
    tmp(09890) := x"0840";
    tmp(09891) := x"0840";
    tmp(09892) := x"0840";
    tmp(09893) := x"0840";
    tmp(09894) := x"0840";
    tmp(09895) := x"0840";
    tmp(09896) := x"0840";
    tmp(09897) := x"0840";
    tmp(09898) := x"0840";
    tmp(09899) := x"0840";
    tmp(09900) := x"0840";
    tmp(09901) := x"0840";
    tmp(09902) := x"0840";
    tmp(09903) := x"0840";
    tmp(09904) := x"0840";
    tmp(09905) := x"0840";
    tmp(09906) := x"0840";
    tmp(09907) := x"0840";
    tmp(09908) := x"0840";
    tmp(09909) := x"0840";
    tmp(09910) := x"0840";
    tmp(09911) := x"0840";
    tmp(09912) := x"0840";
    tmp(09913) := x"0840";
    tmp(09914) := x"0840";
    tmp(09915) := x"0840";
    tmp(09916) := x"0840";
    tmp(09917) := x"0840";
    tmp(09918) := x"0840";
    tmp(09919) := x"0840";
    tmp(09920) := x"0840";
    tmp(09921) := x"0840";
    tmp(09922) := x"0840";
    tmp(09923) := x"0840";
    tmp(09924) := x"0840";
    tmp(09925) := x"0860";
    tmp(09926) := x"0860";
    tmp(09927) := x"0860";
    tmp(09928) := x"0860";
    tmp(09929) := x"0880";
    tmp(09930) := x"0880";
    tmp(09931) := x"0880";
    tmp(09932) := x"0880";
    tmp(09933) := x"0880";
    tmp(09934) := x"0880";
    tmp(09935) := x"0880";
    tmp(09936) := x"0860";
    tmp(09937) := x"0860";
    tmp(09938) := x"0860";
    tmp(09939) := x"0820";
    tmp(09940) := x"0000";
    tmp(09941) := x"0000";
    tmp(09942) := x"0000";
    tmp(09943) := x"0000";
    tmp(09944) := x"0000";
    tmp(09945) := x"0000";
    tmp(09946) := x"0000";
    tmp(09947) := x"0000";
    tmp(09948) := x"0000";
    tmp(09949) := x"0000";
    tmp(09950) := x"0000";
    tmp(09951) := x"0000";
    tmp(09952) := x"0000";
    tmp(09953) := x"0000";
    tmp(09954) := x"0000";
    tmp(09955) := x"0000";
    tmp(09956) := x"0020";
    tmp(09957) := x"1062";
    tmp(09958) := x"0000";
    tmp(09959) := x"0000";
    tmp(09960) := x"0000";
    tmp(09961) := x"0000";
    tmp(09962) := x"0000";
    tmp(09963) := x"0000";
    tmp(09964) := x"0000";
    tmp(09965) := x"0000";
    tmp(09966) := x"0000";
    tmp(09967) := x"0000";
    tmp(09968) := x"0000";
    tmp(09969) := x"0000";
    tmp(09970) := x"0000";
    tmp(09971) := x"0000";
    tmp(09972) := x"0000";
    tmp(09973) := x"0020";
    tmp(09974) := x"0020";
    tmp(09975) := x"0000";
    tmp(09976) := x"0020";
    tmp(09977) := x"0020";
    tmp(09978) := x"0020";
    tmp(09979) := x"0000";
    tmp(09980) := x"0020";
    tmp(09981) := x"0821";
    tmp(09982) := x"0841";
    tmp(09983) := x"0821";
    tmp(09984) := x"0020";
    tmp(09985) := x"0020";
    tmp(09986) := x"0820";
    tmp(09987) := x"1081";
    tmp(09988) := x"3143";
    tmp(09989) := x"2923";
    tmp(09990) := x"20c3";
    tmp(09991) := x"a40e";
    tmp(09992) := x"be33";
    tmp(09993) := x"10c1";
    tmp(09994) := x"0880";
    tmp(09995) := x"08a0";
    tmp(09996) := x"08c0";
    tmp(09997) := x"08c0";
    tmp(09998) := x"08c0";
    tmp(09999) := x"08e0";
    tmp(10000) := x"08e0";
    tmp(10001) := x"08e0";
    tmp(10002) := x"08e0";
    tmp(10003) := x"08e0";
    tmp(10004) := x"08c0";
    tmp(10005) := x"08c0";
    tmp(10006) := x"08c0";
    tmp(10007) := x"08c0";
    tmp(10008) := x"08c0";
    tmp(10009) := x"08c0";
    tmp(10010) := x"08c0";
    tmp(10011) := x"08a0";
    tmp(10012) := x"08a0";
    tmp(10013) := x"08a0";
    tmp(10014) := x"08a0";
    tmp(10015) := x"08a0";
    tmp(10016) := x"0880";
    tmp(10017) := x"0880";
    tmp(10018) := x"0880";
    tmp(10019) := x"0880";
    tmp(10020) := x"0860";
    tmp(10021) := x"0860";
    tmp(10022) := x"0060";
    tmp(10023) := x"0060";
    tmp(10024) := x"0040";
    tmp(10025) := x"0040";
    tmp(10026) := x"0040";
    tmp(10027) := x"0040";
    tmp(10028) := x"0020";
    tmp(10029) := x"0020";
    tmp(10030) := x"0020";
    tmp(10031) := x"0020";
    tmp(10032) := x"0020";
    tmp(10033) := x"0020";
    tmp(10034) := x"0000";
    tmp(10035) := x"0000";
    tmp(10036) := x"0000";
    tmp(10037) := x"ffff";
    tmp(10038) := x"ffff";
    tmp(10039) := x"ffff";
    tmp(10040) := x"ffff";
    tmp(10041) := x"ffff";
    tmp(10042) := x"ffff";
    tmp(10043) := x"ffff";
    tmp(10044) := x"ffff";
    tmp(10045) := x"ffff";
    tmp(10046) := x"ffff";
    tmp(10047) := x"ffff";
    tmp(10048) := x"ffff";
    tmp(10049) := x"ffff";
    tmp(10050) := x"ffff";
    tmp(10051) := x"ffff";
    tmp(10052) := x"ffff";
    tmp(10053) := x"ffff";
    tmp(10054) := x"ffff";
    tmp(10055) := x"ffff";
    tmp(10056) := x"ffff";
    tmp(10057) := x"ffff";
    tmp(10058) := x"ffff";
    tmp(10059) := x"ffff";
    tmp(10060) := x"ffff";
    tmp(10061) := x"ffff";
    tmp(10062) := x"ffff";
    tmp(10063) := x"ffff";
    tmp(10064) := x"ffff";
    tmp(10065) := x"ffff";
    tmp(10066) := x"ffff";
    tmp(10067) := x"ffff";
    tmp(10068) := x"ffff";
    tmp(10069) := x"ffff";
    tmp(10070) := x"ffff";
    tmp(10071) := x"ffff";
    tmp(10072) := x"ffff";
    tmp(10073) := x"ffff";
    tmp(10074) := x"ffff";
    tmp(10075) := x"ffff";
    tmp(10076) := x"ffff";
    tmp(10077) := x"0020";
    tmp(10078) := x"0820";
    tmp(10079) := x"0820";
    tmp(10080) := x"0000";
    tmp(10081) := x"0000";
    tmp(10082) := x"0000";
    tmp(10083) := x"0000";
    tmp(10084) := x"0000";
    tmp(10085) := x"0000";
    tmp(10086) := x"0000";
    tmp(10087) := x"0000";
    tmp(10088) := x"0020";
    tmp(10089) := x"0021";
    tmp(10090) := x"0041";
    tmp(10091) := x"0041";
    tmp(10092) := x"0882";
    tmp(10093) := x"08a3";
    tmp(10094) := x"08c3";
    tmp(10095) := x"08e3";
    tmp(10096) := x"08a2";
    tmp(10097) := x"0881";
    tmp(10098) := x"0861";
    tmp(10099) := x"0841";
    tmp(10100) := x"0040";
    tmp(10101) := x"0020";
    tmp(10102) := x"0020";
    tmp(10103) := x"0020";
    tmp(10104) := x"0820";
    tmp(10105) := x"0820";
    tmp(10106) := x"0820";
    tmp(10107) := x"0820";
    tmp(10108) := x"0820";
    tmp(10109) := x"0820";
    tmp(10110) := x"0820";
    tmp(10111) := x"0820";
    tmp(10112) := x"0820";
    tmp(10113) := x"0820";
    tmp(10114) := x"0820";
    tmp(10115) := x"0820";
    tmp(10116) := x"0820";
    tmp(10117) := x"0820";
    tmp(10118) := x"0820";
    tmp(10119) := x"0820";
    tmp(10120) := x"0820";
    tmp(10121) := x"0820";
    tmp(10122) := x"0820";
    tmp(10123) := x"0820";
    tmp(10124) := x"0820";
    tmp(10125) := x"0840";
    tmp(10126) := x"0820";
    tmp(10127) := x"0820";
    tmp(10128) := x"0840";
    tmp(10129) := x"0840";
    tmp(10130) := x"0840";
    tmp(10131) := x"0840";
    tmp(10132) := x"0820";
    tmp(10133) := x"0840";
    tmp(10134) := x"0840";
    tmp(10135) := x"0840";
    tmp(10136) := x"0840";
    tmp(10137) := x"0840";
    tmp(10138) := x"0840";
    tmp(10139) := x"0840";
    tmp(10140) := x"0840";
    tmp(10141) := x"0840";
    tmp(10142) := x"0840";
    tmp(10143) := x"0840";
    tmp(10144) := x"0840";
    tmp(10145) := x"0840";
    tmp(10146) := x"0840";
    tmp(10147) := x"0840";
    tmp(10148) := x"0840";
    tmp(10149) := x"0840";
    tmp(10150) := x"0840";
    tmp(10151) := x"0840";
    tmp(10152) := x"0840";
    tmp(10153) := x"0840";
    tmp(10154) := x"0840";
    tmp(10155) := x"0840";
    tmp(10156) := x"0840";
    tmp(10157) := x"0840";
    tmp(10158) := x"0840";
    tmp(10159) := x"0840";
    tmp(10160) := x"0840";
    tmp(10161) := x"0840";
    tmp(10162) := x"0840";
    tmp(10163) := x"0840";
    tmp(10164) := x"0860";
    tmp(10165) := x"0860";
    tmp(10166) := x"0860";
    tmp(10167) := x"0860";
    tmp(10168) := x"0860";
    tmp(10169) := x"0860";
    tmp(10170) := x"0860";
    tmp(10171) := x"0860";
    tmp(10172) := x"0880";
    tmp(10173) := x"0860";
    tmp(10174) := x"0860";
    tmp(10175) := x"0860";
    tmp(10176) := x"0860";
    tmp(10177) := x"0860";
    tmp(10178) := x"0860";
    tmp(10179) := x"0020";
    tmp(10180) := x"0000";
    tmp(10181) := x"0000";
    tmp(10182) := x"0000";
    tmp(10183) := x"0000";
    tmp(10184) := x"0000";
    tmp(10185) := x"0000";
    tmp(10186) := x"0000";
    tmp(10187) := x"0000";
    tmp(10188) := x"0000";
    tmp(10189) := x"0000";
    tmp(10190) := x"0000";
    tmp(10191) := x"0000";
    tmp(10192) := x"0000";
    tmp(10193) := x"0000";
    tmp(10194) := x"0000";
    tmp(10195) := x"0020";
    tmp(10196) := x"0020";
    tmp(10197) := x"0000";
    tmp(10198) := x"0862";
    tmp(10199) := x"0841";
    tmp(10200) := x"0000";
    tmp(10201) := x"0000";
    tmp(10202) := x"0000";
    tmp(10203) := x"0000";
    tmp(10204) := x"0020";
    tmp(10205) := x"0000";
    tmp(10206) := x"0000";
    tmp(10207) := x"0000";
    tmp(10208) := x"0000";
    tmp(10209) := x"0000";
    tmp(10210) := x"0000";
    tmp(10211) := x"0000";
    tmp(10212) := x"0000";
    tmp(10213) := x"0020";
    tmp(10214) := x"0020";
    tmp(10215) := x"0020";
    tmp(10216) := x"0000";
    tmp(10217) := x"0821";
    tmp(10218) := x"0020";
    tmp(10219) := x"0020";
    tmp(10220) := x"0020";
    tmp(10221) := x"0020";
    tmp(10222) := x"0821";
    tmp(10223) := x"0841";
    tmp(10224) := x"0821";
    tmp(10225) := x"0020";
    tmp(10226) := x"0821";
    tmp(10227) := x"0841";
    tmp(10228) := x"2923";
    tmp(10229) := x"3163";
    tmp(10230) := x"18a2";
    tmp(10231) := x"4965";
    tmp(10232) := x"ff18";
    tmp(10233) := x"844b";
    tmp(10234) := x"0880";
    tmp(10235) := x"08a0";
    tmp(10236) := x"08c0";
    tmp(10237) := x"08c0";
    tmp(10238) := x"08c0";
    tmp(10239) := x"08e0";
    tmp(10240) := x"08e0";
    tmp(10241) := x"08e0";
    tmp(10242) := x"08c0";
    tmp(10243) := x"08c0";
    tmp(10244) := x"08c0";
    tmp(10245) := x"08e0";
    tmp(10246) := x"08e0";
    tmp(10247) := x"08c0";
    tmp(10248) := x"08c0";
    tmp(10249) := x"08c0";
    tmp(10250) := x"08c0";
    tmp(10251) := x"08c0";
    tmp(10252) := x"08c0";
    tmp(10253) := x"08c0";
    tmp(10254) := x"08a0";
    tmp(10255) := x"08a0";
    tmp(10256) := x"08a0";
    tmp(10257) := x"08a0";
    tmp(10258) := x"08a0";
    tmp(10259) := x"0880";
    tmp(10260) := x"0880";
    tmp(10261) := x"0880";
    tmp(10262) := x"0860";
    tmp(10263) := x"0060";
    tmp(10264) := x"0060";
    tmp(10265) := x"0040";
    tmp(10266) := x"0040";
    tmp(10267) := x"0040";
    tmp(10268) := x"0040";
    tmp(10269) := x"0040";
    tmp(10270) := x"0020";
    tmp(10271) := x"0020";
    tmp(10272) := x"0020";
    tmp(10273) := x"0020";
    tmp(10274) := x"0020";
    tmp(10275) := x"0020";
    tmp(10276) := x"0000";
    tmp(10277) := x"ffff";
    tmp(10278) := x"ffff";
    tmp(10279) := x"ffff";
    tmp(10280) := x"ffff";
    tmp(10281) := x"ffff";
    tmp(10282) := x"ffff";
    tmp(10283) := x"ffff";
    tmp(10284) := x"ffff";
    tmp(10285) := x"ffff";
    tmp(10286) := x"ffff";
    tmp(10287) := x"ffff";
    tmp(10288) := x"ffff";
    tmp(10289) := x"ffff";
    tmp(10290) := x"ffff";
    tmp(10291) := x"ffff";
    tmp(10292) := x"ffff";
    tmp(10293) := x"ffff";
    tmp(10294) := x"ffff";
    tmp(10295) := x"ffff";
    tmp(10296) := x"ffff";
    tmp(10297) := x"ffff";
    tmp(10298) := x"ffff";
    tmp(10299) := x"ffff";
    tmp(10300) := x"ffff";
    tmp(10301) := x"ffff";
    tmp(10302) := x"ffff";
    tmp(10303) := x"ffff";
    tmp(10304) := x"ffff";
    tmp(10305) := x"ffff";
    tmp(10306) := x"ffff";
    tmp(10307) := x"ffff";
    tmp(10308) := x"ffff";
    tmp(10309) := x"ffff";
    tmp(10310) := x"ffff";
    tmp(10311) := x"ffff";
    tmp(10312) := x"ffff";
    tmp(10313) := x"ffff";
    tmp(10314) := x"ffff";
    tmp(10315) := x"ffff";
    tmp(10316) := x"ffff";
    tmp(10317) := x"0020";
    tmp(10318) := x"0020";
    tmp(10319) := x"0820";
    tmp(10320) := x"0000";
    tmp(10321) := x"0021";
    tmp(10322) := x"0021";
    tmp(10323) := x"0021";
    tmp(10324) := x"0021";
    tmp(10325) := x"0020";
    tmp(10326) := x"0020";
    tmp(10327) := x"0000";
    tmp(10328) := x"0000";
    tmp(10329) := x"0000";
    tmp(10330) := x"0000";
    tmp(10331) := x"0020";
    tmp(10332) := x"0021";
    tmp(10333) := x"0021";
    tmp(10334) := x"0041";
    tmp(10335) := x"0883";
    tmp(10336) := x"08e5";
    tmp(10337) := x"0947";
    tmp(10338) := x"1187";
    tmp(10339) := x"0966";
    tmp(10340) := x"0925";
    tmp(10341) := x"08e3";
    tmp(10342) := x"08a2";
    tmp(10343) := x"0861";
    tmp(10344) := x"0841";
    tmp(10345) := x"0820";
    tmp(10346) := x"0020";
    tmp(10347) := x"0820";
    tmp(10348) := x"0820";
    tmp(10349) := x"0820";
    tmp(10350) := x"0820";
    tmp(10351) := x"0820";
    tmp(10352) := x"0820";
    tmp(10353) := x"0820";
    tmp(10354) := x"0820";
    tmp(10355) := x"0820";
    tmp(10356) := x"0820";
    tmp(10357) := x"0820";
    tmp(10358) := x"0820";
    tmp(10359) := x"0820";
    tmp(10360) := x"0820";
    tmp(10361) := x"0820";
    tmp(10362) := x"0820";
    tmp(10363) := x"0820";
    tmp(10364) := x"0820";
    tmp(10365) := x"0820";
    tmp(10366) := x"0820";
    tmp(10367) := x"0820";
    tmp(10368) := x"0820";
    tmp(10369) := x"0820";
    tmp(10370) := x"0840";
    tmp(10371) := x"0820";
    tmp(10372) := x"0840";
    tmp(10373) := x"0840";
    tmp(10374) := x"0820";
    tmp(10375) := x"0840";
    tmp(10376) := x"0840";
    tmp(10377) := x"0840";
    tmp(10378) := x"0840";
    tmp(10379) := x"0840";
    tmp(10380) := x"0840";
    tmp(10381) := x"0840";
    tmp(10382) := x"0840";
    tmp(10383) := x"0840";
    tmp(10384) := x"0840";
    tmp(10385) := x"0840";
    tmp(10386) := x"0840";
    tmp(10387) := x"0840";
    tmp(10388) := x"0840";
    tmp(10389) := x"0840";
    tmp(10390) := x"0840";
    tmp(10391) := x"0840";
    tmp(10392) := x"0840";
    tmp(10393) := x"0840";
    tmp(10394) := x"0840";
    tmp(10395) := x"0840";
    tmp(10396) := x"0840";
    tmp(10397) := x"0840";
    tmp(10398) := x"0840";
    tmp(10399) := x"0840";
    tmp(10400) := x"0840";
    tmp(10401) := x"0840";
    tmp(10402) := x"0840";
    tmp(10403) := x"0840";
    tmp(10404) := x"0840";
    tmp(10405) := x"0860";
    tmp(10406) := x"0860";
    tmp(10407) := x"0860";
    tmp(10408) := x"0860";
    tmp(10409) := x"0860";
    tmp(10410) := x"0840";
    tmp(10411) := x"0840";
    tmp(10412) := x"0860";
    tmp(10413) := x"0860";
    tmp(10414) := x"0860";
    tmp(10415) := x"0860";
    tmp(10416) := x"0860";
    tmp(10417) := x"0860";
    tmp(10418) := x"0860";
    tmp(10419) := x"0020";
    tmp(10420) := x"0000";
    tmp(10421) := x"0000";
    tmp(10422) := x"0000";
    tmp(10423) := x"0000";
    tmp(10424) := x"0000";
    tmp(10425) := x"0000";
    tmp(10426) := x"0000";
    tmp(10427) := x"0000";
    tmp(10428) := x"0000";
    tmp(10429) := x"0000";
    tmp(10430) := x"0000";
    tmp(10431) := x"0000";
    tmp(10432) := x"0000";
    tmp(10433) := x"0000";
    tmp(10434) := x"0000";
    tmp(10435) := x"0000";
    tmp(10436) := x"0020";
    tmp(10437) := x"0020";
    tmp(10438) := x"0000";
    tmp(10439) := x"0841";
    tmp(10440) := x"0861";
    tmp(10441) := x"0000";
    tmp(10442) := x"0000";
    tmp(10443) := x"0000";
    tmp(10444) := x"0000";
    tmp(10445) := x"0000";
    tmp(10446) := x"0000";
    tmp(10447) := x"0000";
    tmp(10448) := x"0020";
    tmp(10449) := x"0000";
    tmp(10450) := x"0000";
    tmp(10451) := x"0000";
    tmp(10452) := x"0020";
    tmp(10453) := x"0020";
    tmp(10454) := x"0000";
    tmp(10455) := x"0020";
    tmp(10456) := x"0020";
    tmp(10457) := x"0020";
    tmp(10458) := x"0821";
    tmp(10459) := x"0020";
    tmp(10460) := x"0000";
    tmp(10461) := x"0020";
    tmp(10462) := x"0841";
    tmp(10463) := x"0841";
    tmp(10464) := x"0821";
    tmp(10465) := x"0020";
    tmp(10466) := x"0821";
    tmp(10467) := x"0841";
    tmp(10468) := x"2902";
    tmp(10469) := x"3963";
    tmp(10470) := x"18a2";
    tmp(10471) := x"4985";
    tmp(10472) := x"fffe";
    tmp(10473) := x"c636";
    tmp(10474) := x"10a1";
    tmp(10475) := x"0860";
    tmp(10476) := x"08a0";
    tmp(10477) := x"08a0";
    tmp(10478) := x"08c0";
    tmp(10479) := x"08c0";
    tmp(10480) := x"08c0";
    tmp(10481) := x"08c0";
    tmp(10482) := x"08c0";
    tmp(10483) := x"08c0";
    tmp(10484) := x"08c0";
    tmp(10485) := x"08c0";
    tmp(10486) := x"08e0";
    tmp(10487) := x"08e0";
    tmp(10488) := x"08e0";
    tmp(10489) := x"08e0";
    tmp(10490) := x"08c0";
    tmp(10491) := x"08c0";
    tmp(10492) := x"08c0";
    tmp(10493) := x"08c0";
    tmp(10494) := x"08c0";
    tmp(10495) := x"08c0";
    tmp(10496) := x"08c0";
    tmp(10497) := x"08a0";
    tmp(10498) := x"08a0";
    tmp(10499) := x"08a0";
    tmp(10500) := x"08a0";
    tmp(10501) := x"08a0";
    tmp(10502) := x"0880";
    tmp(10503) := x"0880";
    tmp(10504) := x"0060";
    tmp(10505) := x"0060";
    tmp(10506) := x"0060";
    tmp(10507) := x"0060";
    tmp(10508) := x"0040";
    tmp(10509) := x"0040";
    tmp(10510) := x"0040";
    tmp(10511) := x"0020";
    tmp(10512) := x"0020";
    tmp(10513) := x"0020";
    tmp(10514) := x"0020";
    tmp(10515) := x"0020";
    tmp(10516) := x"0020";
    tmp(10517) := x"ffff";
    tmp(10518) := x"ffff";
    tmp(10519) := x"ffff";
    tmp(10520) := x"ffff";
    tmp(10521) := x"ffff";
    tmp(10522) := x"ffff";
    tmp(10523) := x"ffff";
    tmp(10524) := x"ffff";
    tmp(10525) := x"ffff";
    tmp(10526) := x"ffff";
    tmp(10527) := x"ffff";
    tmp(10528) := x"ffff";
    tmp(10529) := x"ffff";
    tmp(10530) := x"ffff";
    tmp(10531) := x"ffff";
    tmp(10532) := x"ffff";
    tmp(10533) := x"ffff";
    tmp(10534) := x"ffff";
    tmp(10535) := x"ffff";
    tmp(10536) := x"ffff";
    tmp(10537) := x"ffff";
    tmp(10538) := x"ffff";
    tmp(10539) := x"ffff";
    tmp(10540) := x"ffff";
    tmp(10541) := x"ffff";
    tmp(10542) := x"ffff";
    tmp(10543) := x"ffff";
    tmp(10544) := x"ffff";
    tmp(10545) := x"ffff";
    tmp(10546) := x"ffff";
    tmp(10547) := x"ffff";
    tmp(10548) := x"ffff";
    tmp(10549) := x"ffff";
    tmp(10550) := x"ffff";
    tmp(10551) := x"ffff";
    tmp(10552) := x"ffff";
    tmp(10553) := x"ffff";
    tmp(10554) := x"ffff";
    tmp(10555) := x"ffff";
    tmp(10556) := x"ffff";
    tmp(10557) := x"0020";
    tmp(10558) := x"0020";
    tmp(10559) := x"0820";
    tmp(10560) := x"0000";
    tmp(10561) := x"0085";
    tmp(10562) := x"0065";
    tmp(10563) := x"0065";
    tmp(10564) := x"0064";
    tmp(10565) := x"0064";
    tmp(10566) := x"0063";
    tmp(10567) := x"0043";
    tmp(10568) := x"0042";
    tmp(10569) := x"0041";
    tmp(10570) := x"0021";
    tmp(10571) := x"0021";
    tmp(10572) := x"0021";
    tmp(10573) := x"0021";
    tmp(10574) := x"0021";
    tmp(10575) := x"0041";
    tmp(10576) := x"0082";
    tmp(10577) := x"08c4";
    tmp(10578) := x"08e5";
    tmp(10579) := x"0906";
    tmp(10580) := x"0926";
    tmp(10581) := x"0947";
    tmp(10582) := x"0947";
    tmp(10583) := x"0946";
    tmp(10584) := x"0904";
    tmp(10585) := x"08c3";
    tmp(10586) := x"0882";
    tmp(10587) := x"0861";
    tmp(10588) := x"0861";
    tmp(10589) := x"0841";
    tmp(10590) := x"0820";
    tmp(10591) := x"0820";
    tmp(10592) := x"0820";
    tmp(10593) := x"0820";
    tmp(10594) := x"0820";
    tmp(10595) := x"0820";
    tmp(10596) := x"0820";
    tmp(10597) := x"0820";
    tmp(10598) := x"0820";
    tmp(10599) := x"0820";
    tmp(10600) := x"0820";
    tmp(10601) := x"0820";
    tmp(10602) := x"0820";
    tmp(10603) := x"0820";
    tmp(10604) := x"0820";
    tmp(10605) := x"0820";
    tmp(10606) := x"0820";
    tmp(10607) := x"0820";
    tmp(10608) := x"0820";
    tmp(10609) := x"0820";
    tmp(10610) := x"0820";
    tmp(10611) := x"0820";
    tmp(10612) := x"0820";
    tmp(10613) := x"0820";
    tmp(10614) := x"0820";
    tmp(10615) := x"0820";
    tmp(10616) := x"0820";
    tmp(10617) := x"0840";
    tmp(10618) := x"0840";
    tmp(10619) := x"0840";
    tmp(10620) := x"0840";
    tmp(10621) := x"0840";
    tmp(10622) := x"0840";
    tmp(10623) := x"0840";
    tmp(10624) := x"0840";
    tmp(10625) := x"0840";
    tmp(10626) := x"0840";
    tmp(10627) := x"0840";
    tmp(10628) := x"0840";
    tmp(10629) := x"0840";
    tmp(10630) := x"0840";
    tmp(10631) := x"0840";
    tmp(10632) := x"0840";
    tmp(10633) := x"0840";
    tmp(10634) := x"0840";
    tmp(10635) := x"0840";
    tmp(10636) := x"0840";
    tmp(10637) := x"0840";
    tmp(10638) := x"0840";
    tmp(10639) := x"0840";
    tmp(10640) := x"0840";
    tmp(10641) := x"0840";
    tmp(10642) := x"0840";
    tmp(10643) := x"0840";
    tmp(10644) := x"0840";
    tmp(10645) := x"0860";
    tmp(10646) := x"0840";
    tmp(10647) := x"0840";
    tmp(10648) := x"0820";
    tmp(10649) := x"0840";
    tmp(10650) := x"0840";
    tmp(10651) := x"0820";
    tmp(10652) := x"0820";
    tmp(10653) := x"0840";
    tmp(10654) := x"0840";
    tmp(10655) := x"0860";
    tmp(10656) := x"0860";
    tmp(10657) := x"0860";
    tmp(10658) := x"0840";
    tmp(10659) := x"0000";
    tmp(10660) := x"0000";
    tmp(10661) := x"0000";
    tmp(10662) := x"0000";
    tmp(10663) := x"0000";
    tmp(10664) := x"0000";
    tmp(10665) := x"0000";
    tmp(10666) := x"0000";
    tmp(10667) := x"0000";
    tmp(10668) := x"0000";
    tmp(10669) := x"0000";
    tmp(10670) := x"0000";
    tmp(10671) := x"0000";
    tmp(10672) := x"0000";
    tmp(10673) := x"0000";
    tmp(10674) := x"0000";
    tmp(10675) := x"0000";
    tmp(10676) := x"0000";
    tmp(10677) := x"0000";
    tmp(10678) := x"0000";
    tmp(10679) := x"0020";
    tmp(10680) := x"0841";
    tmp(10681) := x"0000";
    tmp(10682) := x"0000";
    tmp(10683) := x"0000";
    tmp(10684) := x"0000";
    tmp(10685) := x"0000";
    tmp(10686) := x"0000";
    tmp(10687) := x"0000";
    tmp(10688) := x"0020";
    tmp(10689) := x"0020";
    tmp(10690) := x"0000";
    tmp(10691) := x"0020";
    tmp(10692) := x"0020";
    tmp(10693) := x"0020";
    tmp(10694) := x"0000";
    tmp(10695) := x"0020";
    tmp(10696) := x"0020";
    tmp(10697) := x"0000";
    tmp(10698) := x"0020";
    tmp(10699) := x"0020";
    tmp(10700) := x"0020";
    tmp(10701) := x"0020";
    tmp(10702) := x"0821";
    tmp(10703) := x"0841";
    tmp(10704) := x"0841";
    tmp(10705) := x"0821";
    tmp(10706) := x"0821";
    tmp(10707) := x"0841";
    tmp(10708) := x"1881";
    tmp(10709) := x"1881";
    tmp(10710) := x"28e3";
    tmp(10711) := x"8b8c";
    tmp(10712) := x"ffff";
    tmp(10713) := x"c5f4";
    tmp(10714) := x"18c1";
    tmp(10715) := x"08a0";
    tmp(10716) := x"08a0";
    tmp(10717) := x"08a0";
    tmp(10718) := x"08a0";
    tmp(10719) := x"08a0";
    tmp(10720) := x"08c0";
    tmp(10721) := x"08c0";
    tmp(10722) := x"08c0";
    tmp(10723) := x"08c0";
    tmp(10724) := x"08c0";
    tmp(10725) := x"08c0";
    tmp(10726) := x"08c0";
    tmp(10727) := x"08c0";
    tmp(10728) := x"08e0";
    tmp(10729) := x"08c0";
    tmp(10730) := x"08c0";
    tmp(10731) := x"08c0";
    tmp(10732) := x"08c0";
    tmp(10733) := x"08c0";
    tmp(10734) := x"08c0";
    tmp(10735) := x"08c0";
    tmp(10736) := x"08c0";
    tmp(10737) := x"08c0";
    tmp(10738) := x"08c0";
    tmp(10739) := x"08c0";
    tmp(10740) := x"08a0";
    tmp(10741) := x"08a0";
    tmp(10742) := x"08a0";
    tmp(10743) := x"08a0";
    tmp(10744) := x"0880";
    tmp(10745) := x"0880";
    tmp(10746) := x"0060";
    tmp(10747) := x"0060";
    tmp(10748) := x"0060";
    tmp(10749) := x"0060";
    tmp(10750) := x"0040";
    tmp(10751) := x"0040";
    tmp(10752) := x"0040";
    tmp(10753) := x"0040";
    tmp(10754) := x"0020";
    tmp(10755) := x"0020";
    tmp(10756) := x"0020";
    tmp(10757) := x"0000";
    tmp(10758) := x"0000";
    tmp(10759) := x"0000";
    tmp(10760) := x"0000";
    tmp(10761) := x"0000";
    tmp(10762) := x"0000";
    tmp(10763) := x"0000";
    tmp(10764) := x"0000";
    tmp(10765) := x"0000";
    tmp(10766) := x"0000";
    tmp(10767) := x"0000";
    tmp(10768) := x"0000";
    tmp(10769) := x"0000";
    tmp(10770) := x"0000";
    tmp(10771) := x"0000";
    tmp(10772) := x"0000";
    tmp(10773) := x"0000";
    tmp(10774) := x"0000";
    tmp(10775) := x"0000";
    tmp(10776) := x"0000";
    tmp(10777) := x"0000";
    tmp(10778) := x"0000";
    tmp(10779) := x"0000";
    tmp(10780) := x"0000";
    tmp(10781) := x"0000";
    tmp(10782) := x"0000";
    tmp(10783) := x"0000";
    tmp(10784) := x"0000";
    tmp(10785) := x"0000";
    tmp(10786) := x"0000";
    tmp(10787) := x"0000";
    tmp(10788) := x"0000";
    tmp(10789) := x"0000";
    tmp(10790) := x"0000";
    tmp(10791) := x"0000";
    tmp(10792) := x"0000";
    tmp(10793) := x"0000";
    tmp(10794) := x"0000";
    tmp(10795) := x"0000";
    tmp(10796) := x"0000";
    tmp(10797) := x"0020";
    tmp(10798) := x"0020";
    tmp(10799) := x"0820";
    tmp(10800) := x"0000";
    tmp(10801) := x"0043";
    tmp(10802) := x"0063";
    tmp(10803) := x"0063";
    tmp(10804) := x"0063";
    tmp(10805) := x"0064";
    tmp(10806) := x"0064";
    tmp(10807) := x"0064";
    tmp(10808) := x"0065";
    tmp(10809) := x"0065";
    tmp(10810) := x"0064";
    tmp(10811) := x"0064";
    tmp(10812) := x"0062";
    tmp(10813) := x"0882";
    tmp(10814) := x"0882";
    tmp(10815) := x"08a2";
    tmp(10816) := x"0082";
    tmp(10817) := x"0062";
    tmp(10818) := x"0082";
    tmp(10819) := x"0082";
    tmp(10820) := x"0082";
    tmp(10821) := x"0083";
    tmp(10822) := x"00a3";
    tmp(10823) := x"08c4";
    tmp(10824) := x"08e5";
    tmp(10825) := x"0906";
    tmp(10826) := x"0905";
    tmp(10827) := x"08e4";
    tmp(10828) := x"08e4";
    tmp(10829) := x"08c3";
    tmp(10830) := x"08a2";
    tmp(10831) := x"0882";
    tmp(10832) := x"0861";
    tmp(10833) := x"0840";
    tmp(10834) := x"0820";
    tmp(10835) := x"0820";
    tmp(10836) := x"0820";
    tmp(10837) := x"0820";
    tmp(10838) := x"0820";
    tmp(10839) := x"0820";
    tmp(10840) := x"0820";
    tmp(10841) := x"0820";
    tmp(10842) := x"0820";
    tmp(10843) := x"0820";
    tmp(10844) := x"0820";
    tmp(10845) := x"0820";
    tmp(10846) := x"0820";
    tmp(10847) := x"0820";
    tmp(10848) := x"0820";
    tmp(10849) := x"0820";
    tmp(10850) := x"0820";
    tmp(10851) := x"0820";
    tmp(10852) := x"0820";
    tmp(10853) := x"0820";
    tmp(10854) := x"0820";
    tmp(10855) := x"0820";
    tmp(10856) := x"0820";
    tmp(10857) := x"0840";
    tmp(10858) := x"0840";
    tmp(10859) := x"0840";
    tmp(10860) := x"0820";
    tmp(10861) := x"0840";
    tmp(10862) := x"0840";
    tmp(10863) := x"0840";
    tmp(10864) := x"0840";
    tmp(10865) := x"0840";
    tmp(10866) := x"0840";
    tmp(10867) := x"0840";
    tmp(10868) := x"0840";
    tmp(10869) := x"0840";
    tmp(10870) := x"0840";
    tmp(10871) := x"0840";
    tmp(10872) := x"0840";
    tmp(10873) := x"0840";
    tmp(10874) := x"0840";
    tmp(10875) := x"0840";
    tmp(10876) := x"0840";
    tmp(10877) := x"0840";
    tmp(10878) := x"0840";
    tmp(10879) := x"0840";
    tmp(10880) := x"0840";
    tmp(10881) := x"0840";
    tmp(10882) := x"0840";
    tmp(10883) := x"0840";
    tmp(10884) := x"0840";
    tmp(10885) := x"0840";
    tmp(10886) := x"0020";
    tmp(10887) := x"0020";
    tmp(10888) := x"0000";
    tmp(10889) := x"0000";
    tmp(10890) := x"0020";
    tmp(10891) := x"0020";
    tmp(10892) := x"0020";
    tmp(10893) := x"0020";
    tmp(10894) := x"0020";
    tmp(10895) := x"0020";
    tmp(10896) := x"0020";
    tmp(10897) := x"0820";
    tmp(10898) := x"0820";
    tmp(10899) := x"0000";
    tmp(10900) := x"0000";
    tmp(10901) := x"0000";
    tmp(10902) := x"0000";
    tmp(10903) := x"0000";
    tmp(10904) := x"0000";
    tmp(10905) := x"0000";
    tmp(10906) := x"0000";
    tmp(10907) := x"0000";
    tmp(10908) := x"0000";
    tmp(10909) := x"0000";
    tmp(10910) := x"0000";
    tmp(10911) := x"0000";
    tmp(10912) := x"0000";
    tmp(10913) := x"0000";
    tmp(10914) := x"0000";
    tmp(10915) := x"0000";
    tmp(10916) := x"0000";
    tmp(10917) := x"0000";
    tmp(10918) := x"0000";
    tmp(10919) := x"0000";
    tmp(10920) := x"0020";
    tmp(10921) := x"0841";
    tmp(10922) := x"0000";
    tmp(10923) := x"0000";
    tmp(10924) := x"0000";
    tmp(10925) := x"0020";
    tmp(10926) := x"0000";
    tmp(10927) := x"0000";
    tmp(10928) := x"0000";
    tmp(10929) := x"0020";
    tmp(10930) := x"0020";
    tmp(10931) := x"0020";
    tmp(10932) := x"0020";
    tmp(10933) := x"0020";
    tmp(10934) := x"0000";
    tmp(10935) := x"0020";
    tmp(10936) := x"0000";
    tmp(10937) := x"0000";
    tmp(10938) := x"0020";
    tmp(10939) := x"0821";
    tmp(10940) := x"0020";
    tmp(10941) := x"0020";
    tmp(10942) := x"0821";
    tmp(10943) := x"0861";
    tmp(10944) := x"0861";
    tmp(10945) := x"0841";
    tmp(10946) := x"0820";
    tmp(10947) := x"0841";
    tmp(10948) := x"1061";
    tmp(10949) := x"18a2";
    tmp(10950) := x"9c50";
    tmp(10951) := x"ffff";
    tmp(10952) := x"ffff";
    tmp(10953) := x"a4d1";
    tmp(10954) := x"1061";
    tmp(10955) := x"10e1";
    tmp(10956) := x"0880";
    tmp(10957) := x"0880";
    tmp(10958) := x"0880";
    tmp(10959) := x"08a0";
    tmp(10960) := x"08a0";
    tmp(10961) := x"08a0";
    tmp(10962) := x"08a0";
    tmp(10963) := x"08c0";
    tmp(10964) := x"08c0";
    tmp(10965) := x"08c0";
    tmp(10966) := x"08c0";
    tmp(10967) := x"08c0";
    tmp(10968) := x"08c0";
    tmp(10969) := x"08c0";
    tmp(10970) := x"08c0";
    tmp(10971) := x"08c0";
    tmp(10972) := x"08c0";
    tmp(10973) := x"08c0";
    tmp(10974) := x"08c0";
    tmp(10975) := x"08c0";
    tmp(10976) := x"08c0";
    tmp(10977) := x"08c0";
    tmp(10978) := x"08c0";
    tmp(10979) := x"08c0";
    tmp(10980) := x"08c0";
    tmp(10981) := x"08a0";
    tmp(10982) := x"08a0";
    tmp(10983) := x"08a0";
    tmp(10984) := x"08a0";
    tmp(10985) := x"08a0";
    tmp(10986) := x"0880";
    tmp(10987) := x"0880";
    tmp(10988) := x"0080";
    tmp(10989) := x"0060";
    tmp(10990) := x"0060";
    tmp(10991) := x"0060";
    tmp(10992) := x"0040";
    tmp(10993) := x"0040";
    tmp(10994) := x"0040";
    tmp(10995) := x"0020";
    tmp(10996) := x"0020";
    tmp(10997) := x"0000";
    tmp(10998) := x"0000";
    tmp(10999) := x"0000";
    tmp(11000) := x"0000";
    tmp(11001) := x"0000";
    tmp(11002) := x"0000";
    tmp(11003) := x"0000";
    tmp(11004) := x"0000";
    tmp(11005) := x"0000";
    tmp(11006) := x"0000";
    tmp(11007) := x"0000";
    tmp(11008) := x"0000";
    tmp(11009) := x"0000";
    tmp(11010) := x"0000";
    tmp(11011) := x"0000";
    tmp(11012) := x"0000";
    tmp(11013) := x"0000";
    tmp(11014) := x"0000";
    tmp(11015) := x"0000";
    tmp(11016) := x"0000";
    tmp(11017) := x"0000";
    tmp(11018) := x"0000";
    tmp(11019) := x"0000";
    tmp(11020) := x"0000";
    tmp(11021) := x"0000";
    tmp(11022) := x"0000";
    tmp(11023) := x"0000";
    tmp(11024) := x"0000";
    tmp(11025) := x"0000";
    tmp(11026) := x"0000";
    tmp(11027) := x"0000";
    tmp(11028) := x"0000";
    tmp(11029) := x"0000";
    tmp(11030) := x"0000";
    tmp(11031) := x"0000";
    tmp(11032) := x"0000";
    tmp(11033) := x"0000";
    tmp(11034) := x"0000";
    tmp(11035) := x"0000";
    tmp(11036) := x"0000";
    tmp(11037) := x"0020";
    tmp(11038) := x"0020";
    tmp(11039) := x"0020";
    tmp(11040) := x"0000";
    tmp(11041) := x"0861";
    tmp(11042) := x"0862";
    tmp(11043) := x"0882";
    tmp(11044) := x"0882";
    tmp(11045) := x"0862";
    tmp(11046) := x"0862";
    tmp(11047) := x"0862";
    tmp(11048) := x"0862";
    tmp(11049) := x"0862";
    tmp(11050) := x"0863";
    tmp(11051) := x"08a3";
    tmp(11052) := x"08a3";
    tmp(11053) := x"0882";
    tmp(11054) := x"0882";
    tmp(11055) := x"0082";
    tmp(11056) := x"0062";
    tmp(11057) := x"0062";
    tmp(11058) := x"0062";
    tmp(11059) := x"0061";
    tmp(11060) := x"0061";
    tmp(11061) := x"0061";
    tmp(11062) := x"0061";
    tmp(11063) := x"0062";
    tmp(11064) := x"0062";
    tmp(11065) := x"0062";
    tmp(11066) := x"08a2";
    tmp(11067) := x"0882";
    tmp(11068) := x"08a2";
    tmp(11069) := x"08c3";
    tmp(11070) := x"1125";
    tmp(11071) := x"11a7";
    tmp(11072) := x"11a6";
    tmp(11073) := x"1124";
    tmp(11074) := x"08c2";
    tmp(11075) := x"0861";
    tmp(11076) := x"0840";
    tmp(11077) := x"0820";
    tmp(11078) := x"0820";
    tmp(11079) := x"0820";
    tmp(11080) := x"0820";
    tmp(11081) := x"0820";
    tmp(11082) := x"0820";
    tmp(11083) := x"0820";
    tmp(11084) := x"0820";
    tmp(11085) := x"0820";
    tmp(11086) := x"0820";
    tmp(11087) := x"0820";
    tmp(11088) := x"0820";
    tmp(11089) := x"0820";
    tmp(11090) := x"0820";
    tmp(11091) := x"0820";
    tmp(11092) := x"0820";
    tmp(11093) := x"0820";
    tmp(11094) := x"0820";
    tmp(11095) := x"0820";
    tmp(11096) := x"0840";
    tmp(11097) := x"0820";
    tmp(11098) := x"0820";
    tmp(11099) := x"0820";
    tmp(11100) := x"0840";
    tmp(11101) := x"0840";
    tmp(11102) := x"0820";
    tmp(11103) := x"0840";
    tmp(11104) := x"0840";
    tmp(11105) := x"0840";
    tmp(11106) := x"0840";
    tmp(11107) := x"0840";
    tmp(11108) := x"0840";
    tmp(11109) := x"0840";
    tmp(11110) := x"0840";
    tmp(11111) := x"0840";
    tmp(11112) := x"0840";
    tmp(11113) := x"0840";
    tmp(11114) := x"0840";
    tmp(11115) := x"0840";
    tmp(11116) := x"0840";
    tmp(11117) := x"0840";
    tmp(11118) := x"0840";
    tmp(11119) := x"0840";
    tmp(11120) := x"0840";
    tmp(11121) := x"0840";
    tmp(11122) := x"0840";
    tmp(11123) := x"0840";
    tmp(11124) := x"0840";
    tmp(11125) := x"0820";
    tmp(11126) := x"0020";
    tmp(11127) := x"0000";
    tmp(11128) := x"0000";
    tmp(11129) := x"0000";
    tmp(11130) := x"0000";
    tmp(11131) := x"0000";
    tmp(11132) := x"0000";
    tmp(11133) := x"0000";
    tmp(11134) := x"0000";
    tmp(11135) := x"0000";
    tmp(11136) := x"0000";
    tmp(11137) := x"0000";
    tmp(11138) := x"0020";
    tmp(11139) := x"0000";
    tmp(11140) := x"0000";
    tmp(11141) := x"0000";
    tmp(11142) := x"0000";
    tmp(11143) := x"0000";
    tmp(11144) := x"0000";
    tmp(11145) := x"0000";
    tmp(11146) := x"0000";
    tmp(11147) := x"0000";
    tmp(11148) := x"0000";
    tmp(11149) := x"0000";
    tmp(11150) := x"0000";
    tmp(11151) := x"0000";
    tmp(11152) := x"0000";
    tmp(11153) := x"0000";
    tmp(11154) := x"0000";
    tmp(11155) := x"0000";
    tmp(11156) := x"0000";
    tmp(11157) := x"0000";
    tmp(11158) := x"0000";
    tmp(11159) := x"0000";
    tmp(11160) := x"0000";
    tmp(11161) := x"1061";
    tmp(11162) := x"0000";
    tmp(11163) := x"0000";
    tmp(11164) := x"0000";
    tmp(11165) := x"0000";
    tmp(11166) := x"0000";
    tmp(11167) := x"0000";
    tmp(11168) := x"0000";
    tmp(11169) := x"0000";
    tmp(11170) := x"0020";
    tmp(11171) := x"0020";
    tmp(11172) := x"0020";
    tmp(11173) := x"0020";
    tmp(11174) := x"0000";
    tmp(11175) := x"0000";
    tmp(11176) := x"0000";
    tmp(11177) := x"0020";
    tmp(11178) := x"0020";
    tmp(11179) := x"0821";
    tmp(11180) := x"0821";
    tmp(11181) := x"0020";
    tmp(11182) := x"0821";
    tmp(11183) := x"1082";
    tmp(11184) := x"20e4";
    tmp(11185) := x"2925";
    tmp(11186) := x"2904";
    tmp(11187) := x"49e7";
    tmp(11188) := x"836c";
    tmp(11189) := x"ef3b";
    tmp(11190) := x"ffff";
    tmp(11191) := x"ffff";
    tmp(11192) := x"ef7d";
    tmp(11193) := x"49e6";
    tmp(11194) := x"0820";
    tmp(11195) := x"10c1";
    tmp(11196) := x"08c0";
    tmp(11197) := x"0060";
    tmp(11198) := x"0880";
    tmp(11199) := x"0880";
    tmp(11200) := x"0880";
    tmp(11201) := x"0880";
    tmp(11202) := x"08a0";
    tmp(11203) := x"08a0";
    tmp(11204) := x"08a0";
    tmp(11205) := x"08a0";
    tmp(11206) := x"08a0";
    tmp(11207) := x"08c0";
    tmp(11208) := x"08c0";
    tmp(11209) := x"08c0";
    tmp(11210) := x"08c0";
    tmp(11211) := x"08c0";
    tmp(11212) := x"08c0";
    tmp(11213) := x"08c0";
    tmp(11214) := x"08c0";
    tmp(11215) := x"08c0";
    tmp(11216) := x"08c0";
    tmp(11217) := x"08c0";
    tmp(11218) := x"08c0";
    tmp(11219) := x"08c0";
    tmp(11220) := x"08c0";
    tmp(11221) := x"08c0";
    tmp(11222) := x"08c0";
    tmp(11223) := x"08c0";
    tmp(11224) := x"08a0";
    tmp(11225) := x"08a0";
    tmp(11226) := x"08a0";
    tmp(11227) := x"08a0";
    tmp(11228) := x"0880";
    tmp(11229) := x"0080";
    tmp(11230) := x"0080";
    tmp(11231) := x"0060";
    tmp(11232) := x"0060";
    tmp(11233) := x"0060";
    tmp(11234) := x"0040";
    tmp(11235) := x"0040";
    tmp(11236) := x"0040";
    tmp(11237) := x"0000";
    tmp(11238) := x"0000";
    tmp(11239) := x"0000";
    tmp(11240) := x"0000";
    tmp(11241) := x"0000";
    tmp(11242) := x"0000";
    tmp(11243) := x"0000";
    tmp(11244) := x"0000";
    tmp(11245) := x"0000";
    tmp(11246) := x"0000";
    tmp(11247) := x"0000";
    tmp(11248) := x"0000";
    tmp(11249) := x"0000";
    tmp(11250) := x"0000";
    tmp(11251) := x"0000";
    tmp(11252) := x"0000";
    tmp(11253) := x"0000";
    tmp(11254) := x"0000";
    tmp(11255) := x"0000";
    tmp(11256) := x"0000";
    tmp(11257) := x"0000";
    tmp(11258) := x"0000";
    tmp(11259) := x"0000";
    tmp(11260) := x"0000";
    tmp(11261) := x"0000";
    tmp(11262) := x"0000";
    tmp(11263) := x"0000";
    tmp(11264) := x"0000";
    tmp(11265) := x"0000";
    tmp(11266) := x"0000";
    tmp(11267) := x"0000";
    tmp(11268) := x"0000";
    tmp(11269) := x"0000";
    tmp(11270) := x"0000";
    tmp(11271) := x"0000";
    tmp(11272) := x"0000";
    tmp(11273) := x"0000";
    tmp(11274) := x"0000";
    tmp(11275) := x"0000";
    tmp(11276) := x"0000";
    tmp(11277) := x"0020";
    tmp(11278) := x"0020";
    tmp(11279) := x"0020";
    tmp(11280) := x"0000";
    tmp(11281) := x"0841";
    tmp(11282) := x"0841";
    tmp(11283) := x"0841";
    tmp(11284) := x"0841";
    tmp(11285) := x"0841";
    tmp(11286) := x"0841";
    tmp(11287) := x"0861";
    tmp(11288) := x"10a2";
    tmp(11289) := x"18c2";
    tmp(11290) := x"2102";
    tmp(11291) := x"3183";
    tmp(11292) := x"41e3";
    tmp(11293) := x"3a04";
    tmp(11294) := x"2183";
    tmp(11295) := x"08a1";
    tmp(11296) := x"0061";
    tmp(11297) := x"0061";
    tmp(11298) := x"0061";
    tmp(11299) := x"0061";
    tmp(11300) := x"0861";
    tmp(11301) := x"0861";
    tmp(11302) := x"0861";
    tmp(11303) := x"0861";
    tmp(11304) := x"0861";
    tmp(11305) := x"0861";
    tmp(11306) := x"0880";
    tmp(11307) := x"10a0";
    tmp(11308) := x"10a0";
    tmp(11309) := x"10c1";
    tmp(11310) := x"1901";
    tmp(11311) := x"1163";
    tmp(11312) := x"1166";
    tmp(11313) := x"1188";
    tmp(11314) := x"11a8";
    tmp(11315) := x"1187";
    tmp(11316) := x"1124";
    tmp(11317) := x"08a2";
    tmp(11318) := x"0861";
    tmp(11319) := x"0840";
    tmp(11320) := x"0820";
    tmp(11321) := x"0820";
    tmp(11322) := x"0820";
    tmp(11323) := x"0820";
    tmp(11324) := x"0820";
    tmp(11325) := x"0820";
    tmp(11326) := x"0820";
    tmp(11327) := x"0820";
    tmp(11328) := x"0820";
    tmp(11329) := x"0820";
    tmp(11330) := x"0820";
    tmp(11331) := x"0820";
    tmp(11332) := x"0820";
    tmp(11333) := x"0820";
    tmp(11334) := x"0820";
    tmp(11335) := x"0820";
    tmp(11336) := x"0820";
    tmp(11337) := x"0820";
    tmp(11338) := x"0820";
    tmp(11339) := x"0820";
    tmp(11340) := x"0820";
    tmp(11341) := x"0840";
    tmp(11342) := x"0820";
    tmp(11343) := x"0840";
    tmp(11344) := x"0820";
    tmp(11345) := x"0840";
    tmp(11346) := x"0840";
    tmp(11347) := x"0840";
    tmp(11348) := x"0840";
    tmp(11349) := x"0840";
    tmp(11350) := x"0840";
    tmp(11351) := x"0840";
    tmp(11352) := x"0840";
    tmp(11353) := x"0840";
    tmp(11354) := x"0840";
    tmp(11355) := x"0840";
    tmp(11356) := x"0840";
    tmp(11357) := x"0840";
    tmp(11358) := x"0840";
    tmp(11359) := x"0840";
    tmp(11360) := x"0840";
    tmp(11361) := x"0840";
    tmp(11362) := x"0840";
    tmp(11363) := x"0840";
    tmp(11364) := x"0840";
    tmp(11365) := x"0020";
    tmp(11366) := x"0000";
    tmp(11367) := x"0000";
    tmp(11368) := x"0000";
    tmp(11369) := x"0000";
    tmp(11370) := x"0000";
    tmp(11371) := x"0000";
    tmp(11372) := x"0000";
    tmp(11373) := x"0000";
    tmp(11374) := x"0000";
    tmp(11375) := x"0000";
    tmp(11376) := x"0000";
    tmp(11377) := x"0000";
    tmp(11378) := x"0020";
    tmp(11379) := x"0000";
    tmp(11380) := x"0000";
    tmp(11381) := x"0000";
    tmp(11382) := x"0000";
    tmp(11383) := x"0000";
    tmp(11384) := x"0000";
    tmp(11385) := x"0000";
    tmp(11386) := x"0000";
    tmp(11387) := x"0000";
    tmp(11388) := x"0000";
    tmp(11389) := x"0000";
    tmp(11390) := x"0000";
    tmp(11391) := x"0000";
    tmp(11392) := x"0000";
    tmp(11393) := x"0000";
    tmp(11394) := x"0000";
    tmp(11395) := x"0000";
    tmp(11396) := x"0000";
    tmp(11397) := x"0000";
    tmp(11398) := x"0000";
    tmp(11399) := x"0000";
    tmp(11400) := x"0000";
    tmp(11401) := x"0841";
    tmp(11402) := x"0841";
    tmp(11403) := x"0000";
    tmp(11404) := x"0000";
    tmp(11405) := x"0000";
    tmp(11406) := x"0000";
    tmp(11407) := x"0000";
    tmp(11408) := x"0000";
    tmp(11409) := x"0000";
    tmp(11410) := x"0020";
    tmp(11411) := x"0020";
    tmp(11412) := x"0020";
    tmp(11413) := x"0020";
    tmp(11414) := x"0000";
    tmp(11415) := x"0000";
    tmp(11416) := x"0000";
    tmp(11417) := x"0000";
    tmp(11418) := x"0020";
    tmp(11419) := x"0020";
    tmp(11420) := x"0020";
    tmp(11421) := x"0841";
    tmp(11422) := x"18c3";
    tmp(11423) := x"49e8";
    tmp(11424) := x"72ed";
    tmp(11425) := x"8b8f";
    tmp(11426) := x"cd55";
    tmp(11427) := x"ffdf";
    tmp(11428) := x"ff1c";
    tmp(11429) := x"ff3c";
    tmp(11430) := x"ff9d";
    tmp(11431) := x"fe98";
    tmp(11432) := x"e636";
    tmp(11433) := x"49e5";
    tmp(11434) := x"0820";
    tmp(11435) := x"0880";
    tmp(11436) := x"1100";
    tmp(11437) := x"0880";
    tmp(11438) := x"0860";
    tmp(11439) := x"0860";
    tmp(11440) := x"0860";
    tmp(11441) := x"0880";
    tmp(11442) := x"0880";
    tmp(11443) := x"0880";
    tmp(11444) := x"0880";
    tmp(11445) := x"0880";
    tmp(11446) := x"08a0";
    tmp(11447) := x"08a0";
    tmp(11448) := x"08a0";
    tmp(11449) := x"08a0";
    tmp(11450) := x"08a0";
    tmp(11451) := x"08a0";
    tmp(11452) := x"08c0";
    tmp(11453) := x"08c0";
    tmp(11454) := x"08c0";
    tmp(11455) := x"08c0";
    tmp(11456) := x"08c0";
    tmp(11457) := x"08c0";
    tmp(11458) := x"08c0";
    tmp(11459) := x"08c0";
    tmp(11460) := x"08c0";
    tmp(11461) := x"08c0";
    tmp(11462) := x"08c0";
    tmp(11463) := x"08c0";
    tmp(11464) := x"08a0";
    tmp(11465) := x"08a0";
    tmp(11466) := x"08a0";
    tmp(11467) := x"08a0";
    tmp(11468) := x"08a0";
    tmp(11469) := x"0080";
    tmp(11470) := x"0080";
    tmp(11471) := x"0080";
    tmp(11472) := x"0080";
    tmp(11473) := x"0060";
    tmp(11474) := x"0060";
    tmp(11475) := x"0060";
    tmp(11476) := x"0040";
    tmp(11477) := x"0000";
    tmp(11478) := x"0000";
    tmp(11479) := x"0000";
    tmp(11480) := x"0000";
    tmp(11481) := x"0000";
    tmp(11482) := x"0000";
    tmp(11483) := x"0000";
    tmp(11484) := x"0000";
    tmp(11485) := x"0000";
    tmp(11486) := x"0000";
    tmp(11487) := x"0000";
    tmp(11488) := x"0000";
    tmp(11489) := x"0000";
    tmp(11490) := x"0000";
    tmp(11491) := x"0000";
    tmp(11492) := x"0000";
    tmp(11493) := x"0000";
    tmp(11494) := x"0000";
    tmp(11495) := x"0000";
    tmp(11496) := x"0000";
    tmp(11497) := x"0000";
    tmp(11498) := x"0000";
    tmp(11499) := x"0000";
    tmp(11500) := x"0000";
    tmp(11501) := x"0000";
    tmp(11502) := x"0000";
    tmp(11503) := x"0000";
    tmp(11504) := x"0000";
    tmp(11505) := x"0000";
    tmp(11506) := x"0000";
    tmp(11507) := x"0000";
    tmp(11508) := x"0000";
    tmp(11509) := x"0000";
    tmp(11510) := x"0000";
    tmp(11511) := x"0000";
    tmp(11512) := x"0000";
    tmp(11513) := x"0000";
    tmp(11514) := x"0000";
    tmp(11515) := x"0000";
    tmp(11516) := x"0000";
    tmp(11517) := x"0020";
    tmp(11518) := x"0020";
    tmp(11519) := x"0020";
    tmp(11520) := x"0000";
    tmp(11521) := x"0041";
    tmp(11522) := x"0020";
    tmp(11523) := x"0020";
    tmp(11524) := x"0020";
    tmp(11525) := x"0020";
    tmp(11526) := x"0020";
    tmp(11527) := x"0841";
    tmp(11528) := x"0861";
    tmp(11529) := x"1081";
    tmp(11530) := x"20c1";
    tmp(11531) := x"3142";
    tmp(11532) := x"51e2";
    tmp(11533) := x"6283";
    tmp(11534) := x"7304";
    tmp(11535) := x"4a22";
    tmp(11536) := x"2101";
    tmp(11537) := x"10a0";
    tmp(11538) := x"10a0";
    tmp(11539) := x"10a0";
    tmp(11540) := x"10a0";
    tmp(11541) := x"18c0";
    tmp(11542) := x"18c0";
    tmp(11543) := x"18a0";
    tmp(11544) := x"18c0";
    tmp(11545) := x"20e0";
    tmp(11546) := x"20e0";
    tmp(11547) := x"2900";
    tmp(11548) := x"2900";
    tmp(11549) := x"2900";
    tmp(11550) := x"2920";
    tmp(11551) := x"2920";
    tmp(11552) := x"1921";
    tmp(11553) := x"1102";
    tmp(11554) := x"08e3";
    tmp(11555) := x"1146";
    tmp(11556) := x"1187";
    tmp(11557) := x"11a7";
    tmp(11558) := x"1186";
    tmp(11559) := x"1124";
    tmp(11560) := x"08a2";
    tmp(11561) := x"0841";
    tmp(11562) := x"0820";
    tmp(11563) := x"0820";
    tmp(11564) := x"0820";
    tmp(11565) := x"0820";
    tmp(11566) := x"0820";
    tmp(11567) := x"0820";
    tmp(11568) := x"0820";
    tmp(11569) := x"0820";
    tmp(11570) := x"0820";
    tmp(11571) := x"0820";
    tmp(11572) := x"0820";
    tmp(11573) := x"0820";
    tmp(11574) := x"0820";
    tmp(11575) := x"0820";
    tmp(11576) := x"0820";
    tmp(11577) := x"0820";
    tmp(11578) := x"0820";
    tmp(11579) := x"0820";
    tmp(11580) := x"0840";
    tmp(11581) := x"0820";
    tmp(11582) := x"0840";
    tmp(11583) := x"0820";
    tmp(11584) := x"0820";
    tmp(11585) := x"0820";
    tmp(11586) := x"0820";
    tmp(11587) := x"0820";
    tmp(11588) := x"0820";
    tmp(11589) := x"0820";
    tmp(11590) := x"0820";
    tmp(11591) := x"0840";
    tmp(11592) := x"0820";
    tmp(11593) := x"0840";
    tmp(11594) := x"0840";
    tmp(11595) := x"0840";
    tmp(11596) := x"0840";
    tmp(11597) := x"0840";
    tmp(11598) := x"0840";
    tmp(11599) := x"0840";
    tmp(11600) := x"0840";
    tmp(11601) := x"0840";
    tmp(11602) := x"0840";
    tmp(11603) := x"0840";
    tmp(11604) := x"0020";
    tmp(11605) := x"0000";
    tmp(11606) := x"0000";
    tmp(11607) := x"0000";
    tmp(11608) := x"0000";
    tmp(11609) := x"0000";
    tmp(11610) := x"0000";
    tmp(11611) := x"0000";
    tmp(11612) := x"0000";
    tmp(11613) := x"0000";
    tmp(11614) := x"0000";
    tmp(11615) := x"0000";
    tmp(11616) := x"0000";
    tmp(11617) := x"0000";
    tmp(11618) := x"0020";
    tmp(11619) := x"0000";
    tmp(11620) := x"0000";
    tmp(11621) := x"0000";
    tmp(11622) := x"0000";
    tmp(11623) := x"0000";
    tmp(11624) := x"0000";
    tmp(11625) := x"0000";
    tmp(11626) := x"0000";
    tmp(11627) := x"0000";
    tmp(11628) := x"0000";
    tmp(11629) := x"0000";
    tmp(11630) := x"0000";
    tmp(11631) := x"0000";
    tmp(11632) := x"0000";
    tmp(11633) := x"0000";
    tmp(11634) := x"0000";
    tmp(11635) := x"0000";
    tmp(11636) := x"0000";
    tmp(11637) := x"0000";
    tmp(11638) := x"0000";
    tmp(11639) := x"0000";
    tmp(11640) := x"0000";
    tmp(11641) := x"0821";
    tmp(11642) := x"0841";
    tmp(11643) := x"0000";
    tmp(11644) := x"0000";
    tmp(11645) := x"0020";
    tmp(11646) := x"0000";
    tmp(11647) := x"0000";
    tmp(11648) := x"0000";
    tmp(11649) := x"0000";
    tmp(11650) := x"0020";
    tmp(11651) := x"0000";
    tmp(11652) := x"0020";
    tmp(11653) := x"0000";
    tmp(11654) := x"0000";
    tmp(11655) := x"0000";
    tmp(11656) := x"0000";
    tmp(11657) := x"0000";
    tmp(11658) := x"0820";
    tmp(11659) := x"18a2";
    tmp(11660) := x"3145";
    tmp(11661) := x"5249";
    tmp(11662) := x"6acd";
    tmp(11663) := x"8b70";
    tmp(11664) := x"c4d6";
    tmp(11665) := x"b433";
    tmp(11666) := x"cd36";
    tmp(11667) := x"dd77";
    tmp(11668) := x"d493";
    tmp(11669) := x"ed76";
    tmp(11670) := x"fe99";
    tmp(11671) := x"fe97";
    tmp(11672) := x"d531";
    tmp(11673) := x"2903";
    tmp(11674) := x"0840";
    tmp(11675) := x"0860";
    tmp(11676) := x"1920";
    tmp(11677) := x"08a0";
    tmp(11678) := x"0060";
    tmp(11679) := x"0860";
    tmp(11680) := x"0060";
    tmp(11681) := x"0860";
    tmp(11682) := x"0060";
    tmp(11683) := x"0860";
    tmp(11684) := x"0060";
    tmp(11685) := x"0880";
    tmp(11686) := x"0080";
    tmp(11687) := x"0880";
    tmp(11688) := x"0880";
    tmp(11689) := x"0880";
    tmp(11690) := x"08a0";
    tmp(11691) := x"08a0";
    tmp(11692) := x"08a0";
    tmp(11693) := x"08a0";
    tmp(11694) := x"08a0";
    tmp(11695) := x"08a0";
    tmp(11696) := x"08a0";
    tmp(11697) := x"08c0";
    tmp(11698) := x"08c0";
    tmp(11699) := x"08c0";
    tmp(11700) := x"08c0";
    tmp(11701) := x"08c0";
    tmp(11702) := x"08c0";
    tmp(11703) := x"08a0";
    tmp(11704) := x"08a0";
    tmp(11705) := x"08a0";
    tmp(11706) := x"08a0";
    tmp(11707) := x"08a0";
    tmp(11708) := x"08a0";
    tmp(11709) := x"08a0";
    tmp(11710) := x"00a0";
    tmp(11711) := x"0080";
    tmp(11712) := x"0080";
    tmp(11713) := x"0080";
    tmp(11714) := x"0080";
    tmp(11715) := x"0060";
    tmp(11716) := x"0060";
    tmp(11717) := x"0000";
    tmp(11718) := x"0000";
    tmp(11719) := x"0000";
    tmp(11720) := x"0000";
    tmp(11721) := x"0000";
    tmp(11722) := x"0000";
    tmp(11723) := x"0000";
    tmp(11724) := x"0000";
    tmp(11725) := x"0000";
    tmp(11726) := x"0000";
    tmp(11727) := x"0000";
    tmp(11728) := x"0000";
    tmp(11729) := x"0000";
    tmp(11730) := x"0000";
    tmp(11731) := x"0000";
    tmp(11732) := x"0000";
    tmp(11733) := x"0000";
    tmp(11734) := x"0000";
    tmp(11735) := x"0000";
    tmp(11736) := x"0000";
    tmp(11737) := x"0000";
    tmp(11738) := x"0000";
    tmp(11739) := x"0000";
    tmp(11740) := x"0000";
    tmp(11741) := x"0000";
    tmp(11742) := x"0000";
    tmp(11743) := x"0000";
    tmp(11744) := x"0000";
    tmp(11745) := x"0000";
    tmp(11746) := x"0000";
    tmp(11747) := x"0000";
    tmp(11748) := x"0000";
    tmp(11749) := x"0000";
    tmp(11750) := x"0000";
    tmp(11751) := x"0000";
    tmp(11752) := x"0000";
    tmp(11753) := x"0000";
    tmp(11754) := x"0000";
    tmp(11755) := x"0000";
    tmp(11756) := x"0000";
    tmp(11757) := x"0000";
    tmp(11758) := x"0020";
    tmp(11759) := x"0020";
    tmp(11760) := x"0000";
    tmp(11761) := x"0041";
    tmp(11762) := x"0041";
    tmp(11763) := x"0041";
    tmp(11764) := x"0021";
    tmp(11765) := x"0021";
    tmp(11766) := x"0021";
    tmp(11767) := x"0041";
    tmp(11768) := x"0841";
    tmp(11769) := x"1081";
    tmp(11770) := x"18c1";
    tmp(11771) := x"3141";
    tmp(11772) := x"41a1";
    tmp(11773) := x"5a41";
    tmp(11774) := x"7aa1";
    tmp(11775) := x"7aa0";
    tmp(11776) := x"6200";
    tmp(11777) := x"49a0";
    tmp(11778) := x"3940";
    tmp(11779) := x"3120";
    tmp(11780) := x"28e0";
    tmp(11781) := x"3120";
    tmp(11782) := x"3940";
    tmp(11783) := x"4140";
    tmp(11784) := x"3940";
    tmp(11785) := x"3920";
    tmp(11786) := x"4140";
    tmp(11787) := x"4980";
    tmp(11788) := x"5180";
    tmp(11789) := x"4960";
    tmp(11790) := x"5180";
    tmp(11791) := x"4960";
    tmp(11792) := x"4160";
    tmp(11793) := x"3960";
    tmp(11794) := x"2101";
    tmp(11795) := x"1901";
    tmp(11796) := x"2163";
    tmp(11797) := x"1944";
    tmp(11798) := x"1186";
    tmp(11799) := x"19c8";
    tmp(11800) := x"2208";
    tmp(11801) := x"1165";
    tmp(11802) := x"10c2";
    tmp(11803) := x"0861";
    tmp(11804) := x"0840";
    tmp(11805) := x"0840";
    tmp(11806) := x"0840";
    tmp(11807) := x"0820";
    tmp(11808) := x"0820";
    tmp(11809) := x"0820";
    tmp(11810) := x"0820";
    tmp(11811) := x"0820";
    tmp(11812) := x"0820";
    tmp(11813) := x"0820";
    tmp(11814) := x"0820";
    tmp(11815) := x"0820";
    tmp(11816) := x"0820";
    tmp(11817) := x"0820";
    tmp(11818) := x"0820";
    tmp(11819) := x"0820";
    tmp(11820) := x"0820";
    tmp(11821) := x"0820";
    tmp(11822) := x"0820";
    tmp(11823) := x"0820";
    tmp(11824) := x"0820";
    tmp(11825) := x"0820";
    tmp(11826) := x"0820";
    tmp(11827) := x"0820";
    tmp(11828) := x"0820";
    tmp(11829) := x"0820";
    tmp(11830) := x"0840";
    tmp(11831) := x"0820";
    tmp(11832) := x"0820";
    tmp(11833) := x"0840";
    tmp(11834) := x"0840";
    tmp(11835) := x"0840";
    tmp(11836) := x"0840";
    tmp(11837) := x"0840";
    tmp(11838) := x"0840";
    tmp(11839) := x"0840";
    tmp(11840) := x"0840";
    tmp(11841) := x"0840";
    tmp(11842) := x"0840";
    tmp(11843) := x"0020";
    tmp(11844) := x"0000";
    tmp(11845) := x"0000";
    tmp(11846) := x"0000";
    tmp(11847) := x"0000";
    tmp(11848) := x"0000";
    tmp(11849) := x"0000";
    tmp(11850) := x"0000";
    tmp(11851) := x"0000";
    tmp(11852) := x"0000";
    tmp(11853) := x"0000";
    tmp(11854) := x"0000";
    tmp(11855) := x"0000";
    tmp(11856) := x"0000";
    tmp(11857) := x"0020";
    tmp(11858) := x"0841";
    tmp(11859) := x"0000";
    tmp(11860) := x"0000";
    tmp(11861) := x"0000";
    tmp(11862) := x"0000";
    tmp(11863) := x"0000";
    tmp(11864) := x"0000";
    tmp(11865) := x"0000";
    tmp(11866) := x"0000";
    tmp(11867) := x"0000";
    tmp(11868) := x"0000";
    tmp(11869) := x"0000";
    tmp(11870) := x"0000";
    tmp(11871) := x"0000";
    tmp(11872) := x"0000";
    tmp(11873) := x"0000";
    tmp(11874) := x"0000";
    tmp(11875) := x"0000";
    tmp(11876) := x"0000";
    tmp(11877) := x"0000";
    tmp(11878) := x"0000";
    tmp(11879) := x"0000";
    tmp(11880) := x"0000";
    tmp(11881) := x"0020";
    tmp(11882) := x"0841";
    tmp(11883) := x"0020";
    tmp(11884) := x"0820";
    tmp(11885) := x"1082";
    tmp(11886) := x"1061";
    tmp(11887) := x"0020";
    tmp(11888) := x"0000";
    tmp(11889) := x"0020";
    tmp(11890) := x"0000";
    tmp(11891) := x"0000";
    tmp(11892) := x"0000";
    tmp(11893) := x"0000";
    tmp(11894) := x"0000";
    tmp(11895) := x"0000";
    tmp(11896) := x"0841";
    tmp(11897) := x"2904";
    tmp(11898) := x"5208";
    tmp(11899) := x"730d";
    tmp(11900) := x"93b0";
    tmp(11901) := x"93b1";
    tmp(11902) := x"8b50";
    tmp(11903) := x"a3b1";
    tmp(11904) := x"d4d6";
    tmp(11905) := x"c453";
    tmp(11906) := x"c412";
    tmp(11907) := x"cc32";
    tmp(11908) := x"bbb0";
    tmp(11909) := x"e5b7";
    tmp(11910) := x"e4d2";
    tmp(11911) := x"b3ee";
    tmp(11912) := x"7b0a";
    tmp(11913) := x"0820";
    tmp(11914) := x"0860";
    tmp(11915) := x"0860";
    tmp(11916) := x"1921";
    tmp(11917) := x"10e0";
    tmp(11918) := x"0040";
    tmp(11919) := x"0860";
    tmp(11920) := x"0060";
    tmp(11921) := x"0060";
    tmp(11922) := x"0060";
    tmp(11923) := x"0060";
    tmp(11924) := x"0060";
    tmp(11925) := x"0060";
    tmp(11926) := x"0060";
    tmp(11927) := x"0060";
    tmp(11928) := x"0060";
    tmp(11929) := x"0060";
    tmp(11930) := x"0080";
    tmp(11931) := x"0080";
    tmp(11932) := x"0880";
    tmp(11933) := x"0880";
    tmp(11934) := x"08a0";
    tmp(11935) := x"08a0";
    tmp(11936) := x"08a0";
    tmp(11937) := x"08a0";
    tmp(11938) := x"08a0";
    tmp(11939) := x"08a0";
    tmp(11940) := x"08a0";
    tmp(11941) := x"08c0";
    tmp(11942) := x"08c0";
    tmp(11943) := x"08c0";
    tmp(11944) := x"08a0";
    tmp(11945) := x"08a0";
    tmp(11946) := x"08a0";
    tmp(11947) := x"08a0";
    tmp(11948) := x"08a0";
    tmp(11949) := x"08a0";
    tmp(11950) := x"08a0";
    tmp(11951) := x"08a0";
    tmp(11952) := x"0080";
    tmp(11953) := x"0080";
    tmp(11954) := x"0080";
    tmp(11955) := x"0060";
    tmp(11956) := x"0060";
    tmp(11957) := x"0000";
    tmp(11958) := x"0000";
    tmp(11959) := x"0000";
    tmp(11960) := x"0000";
    tmp(11961) := x"0000";
    tmp(11962) := x"0000";
    tmp(11963) := x"0000";
    tmp(11964) := x"0000";
    tmp(11965) := x"0000";
    tmp(11966) := x"0000";
    tmp(11967) := x"0000";
    tmp(11968) := x"0000";
    tmp(11969) := x"0000";
    tmp(11970) := x"0000";
    tmp(11971) := x"0000";
    tmp(11972) := x"0000";
    tmp(11973) := x"0000";
    tmp(11974) := x"0000";
    tmp(11975) := x"0000";
    tmp(11976) := x"0000";
    tmp(11977) := x"0000";
    tmp(11978) := x"0000";
    tmp(11979) := x"0000";
    tmp(11980) := x"0000";
    tmp(11981) := x"0000";
    tmp(11982) := x"0000";
    tmp(11983) := x"0000";
    tmp(11984) := x"0000";
    tmp(11985) := x"0000";
    tmp(11986) := x"0000";
    tmp(11987) := x"0000";
    tmp(11988) := x"0000";
    tmp(11989) := x"0000";
    tmp(11990) := x"0000";
    tmp(11991) := x"0000";
    tmp(11992) := x"0000";
    tmp(11993) := x"0000";
    tmp(11994) := x"0000";
    tmp(11995) := x"0000";
    tmp(11996) := x"0000";
    tmp(11997) := x"0000";
    tmp(11998) := x"0020";
    tmp(11999) := x"0020";
    tmp(12000) := x"0000";
    tmp(12001) := x"0041";
    tmp(12002) := x"0061";
    tmp(12003) := x"0061";
    tmp(12004) := x"0041";
    tmp(12005) := x"0041";
    tmp(12006) := x"0041";
    tmp(12007) := x"0041";
    tmp(12008) := x"0861";
    tmp(12009) := x"0881";
    tmp(12010) := x"18c1";
    tmp(12011) := x"3141";
    tmp(12012) := x"4180";
    tmp(12013) := x"51c0";
    tmp(12014) := x"6200";
    tmp(12015) := x"6a20";
    tmp(12016) := x"6a00";
    tmp(12017) := x"69e0";
    tmp(12018) := x"61c0";
    tmp(12019) := x"59c0";
    tmp(12020) := x"5180";
    tmp(12021) := x"5180";
    tmp(12022) := x"59a0";
    tmp(12023) := x"61c0";
    tmp(12024) := x"59a0";
    tmp(12025) := x"59a0";
    tmp(12026) := x"61a0";
    tmp(12027) := x"61a0";
    tmp(12028) := x"69c0";
    tmp(12029) := x"69a0";
    tmp(12030) := x"61a0";
    tmp(12031) := x"69e0";
    tmp(12032) := x"69c0";
    tmp(12033) := x"6a00";
    tmp(12034) := x"61e0";
    tmp(12035) := x"51c0";
    tmp(12036) := x"51c1";
    tmp(12037) := x"3141";
    tmp(12038) := x"2142";
    tmp(12039) := x"2983";
    tmp(12040) := x"3225";
    tmp(12041) := x"3a87";
    tmp(12042) := x"3205";
    tmp(12043) := x"39c4";
    tmp(12044) := x"39a1";
    tmp(12045) := x"4981";
    tmp(12046) := x"3100";
    tmp(12047) := x"1080";
    tmp(12048) := x"0840";
    tmp(12049) := x"0820";
    tmp(12050) := x"0820";
    tmp(12051) := x"0820";
    tmp(12052) := x"0820";
    tmp(12053) := x"0820";
    tmp(12054) := x"0820";
    tmp(12055) := x"0820";
    tmp(12056) := x"0820";
    tmp(12057) := x"0820";
    tmp(12058) := x"0820";
    tmp(12059) := x"0820";
    tmp(12060) := x"0820";
    tmp(12061) := x"0820";
    tmp(12062) := x"0820";
    tmp(12063) := x"0820";
    tmp(12064) := x"0820";
    tmp(12065) := x"0820";
    tmp(12066) := x"0820";
    tmp(12067) := x"0820";
    tmp(12068) := x"0820";
    tmp(12069) := x"0820";
    tmp(12070) := x"0820";
    tmp(12071) := x"0820";
    tmp(12072) := x"0820";
    tmp(12073) := x"0820";
    tmp(12074) := x"0820";
    tmp(12075) := x"0820";
    tmp(12076) := x"0840";
    tmp(12077) := x"0840";
    tmp(12078) := x"0840";
    tmp(12079) := x"0860";
    tmp(12080) := x"0860";
    tmp(12081) := x"0860";
    tmp(12082) := x"0840";
    tmp(12083) := x"0020";
    tmp(12084) := x"0000";
    tmp(12085) := x"0000";
    tmp(12086) := x"0000";
    tmp(12087) := x"0000";
    tmp(12088) := x"0000";
    tmp(12089) := x"0000";
    tmp(12090) := x"0000";
    tmp(12091) := x"0000";
    tmp(12092) := x"0000";
    tmp(12093) := x"0000";
    tmp(12094) := x"0000";
    tmp(12095) := x"0000";
    tmp(12096) := x"0000";
    tmp(12097) := x"0000";
    tmp(12098) := x"1081";
    tmp(12099) := x"0820";
    tmp(12100) := x"0000";
    tmp(12101) := x"0000";
    tmp(12102) := x"0000";
    tmp(12103) := x"0000";
    tmp(12104) := x"0000";
    tmp(12105) := x"0000";
    tmp(12106) := x"0000";
    tmp(12107) := x"0000";
    tmp(12108) := x"0000";
    tmp(12109) := x"0000";
    tmp(12110) := x"0000";
    tmp(12111) := x"0000";
    tmp(12112) := x"0000";
    tmp(12113) := x"0000";
    tmp(12114) := x"0000";
    tmp(12115) := x"0000";
    tmp(12116) := x"0000";
    tmp(12117) := x"0000";
    tmp(12118) := x"0000";
    tmp(12119) := x"0000";
    tmp(12120) := x"0000";
    tmp(12121) := x"0000";
    tmp(12122) := x"1061";
    tmp(12123) := x"1061";
    tmp(12124) := x"3124";
    tmp(12125) := x"72eb";
    tmp(12126) := x"5a49";
    tmp(12127) := x"3985";
    tmp(12128) := x"20e3";
    tmp(12129) := x"2904";
    tmp(12130) := x"20c3";
    tmp(12131) := x"18a2";
    tmp(12132) := x"20e3";
    tmp(12133) := x"3165";
    tmp(12134) := x"49e7";
    tmp(12135) := x"5208";
    tmp(12136) := x"834d";
    tmp(12137) := x"93b0";
    tmp(12138) := x"ac53";
    tmp(12139) := x"8b70";
    tmp(12140) := x"832f";
    tmp(12141) := x"830e";
    tmp(12142) := x"9b90";
    tmp(12143) := x"cc73";
    tmp(12144) := x"bc11";
    tmp(12145) := x"bbd1";
    tmp(12146) := x"ab4f";
    tmp(12147) := x"8a8b";
    tmp(12148) := x"ab4e";
    tmp(12149) := x"dcf5";
    tmp(12150) := x"e4f2";
    tmp(12151) := x"ab8c";
    tmp(12152) := x"1061";
    tmp(12153) := x"0840";
    tmp(12154) := x"0840";
    tmp(12155) := x"0820";
    tmp(12156) := x"1921";
    tmp(12157) := x"1120";
    tmp(12158) := x"0060";
    tmp(12159) := x"0860";
    tmp(12160) := x"0060";
    tmp(12161) := x"0860";
    tmp(12162) := x"0860";
    tmp(12163) := x"0040";
    tmp(12164) := x"0040";
    tmp(12165) := x"0040";
    tmp(12166) := x"0040";
    tmp(12167) := x"0040";
    tmp(12168) := x"0060";
    tmp(12169) := x"0060";
    tmp(12170) := x"0060";
    tmp(12171) := x"0060";
    tmp(12172) := x"0060";
    tmp(12173) := x"0080";
    tmp(12174) := x"0080";
    tmp(12175) := x"0880";
    tmp(12176) := x"0880";
    tmp(12177) := x"0880";
    tmp(12178) := x"08a0";
    tmp(12179) := x"08a0";
    tmp(12180) := x"08a0";
    tmp(12181) := x"08a0";
    tmp(12182) := x"08a0";
    tmp(12183) := x"08a0";
    tmp(12184) := x"08a0";
    tmp(12185) := x"08a0";
    tmp(12186) := x"08a0";
    tmp(12187) := x"08a0";
    tmp(12188) := x"08a0";
    tmp(12189) := x"08a0";
    tmp(12190) := x"08a0";
    tmp(12191) := x"08a0";
    tmp(12192) := x"0080";
    tmp(12193) := x"0080";
    tmp(12194) := x"0080";
    tmp(12195) := x"0080";
    tmp(12196) := x"0060";
    tmp(12197) := x"0000";
    tmp(12198) := x"0000";
    tmp(12199) := x"0000";
    tmp(12200) := x"0000";
    tmp(12201) := x"0000";
    tmp(12202) := x"0000";
    tmp(12203) := x"0000";
    tmp(12204) := x"0000";
    tmp(12205) := x"0000";
    tmp(12206) := x"0000";
    tmp(12207) := x"0000";
    tmp(12208) := x"0000";
    tmp(12209) := x"0000";
    tmp(12210) := x"0000";
    tmp(12211) := x"0000";
    tmp(12212) := x"0000";
    tmp(12213) := x"0000";
    tmp(12214) := x"0000";
    tmp(12215) := x"0000";
    tmp(12216) := x"0000";
    tmp(12217) := x"0000";
    tmp(12218) := x"0000";
    tmp(12219) := x"0000";
    tmp(12220) := x"0000";
    tmp(12221) := x"0000";
    tmp(12222) := x"0000";
    tmp(12223) := x"0000";
    tmp(12224) := x"0000";
    tmp(12225) := x"0000";
    tmp(12226) := x"0000";
    tmp(12227) := x"0000";
    tmp(12228) := x"0000";
    tmp(12229) := x"0000";
    tmp(12230) := x"0000";
    tmp(12231) := x"0000";
    tmp(12232) := x"0000";
    tmp(12233) := x"0000";
    tmp(12234) := x"0000";
    tmp(12235) := x"0000";
    tmp(12236) := x"0000";
    tmp(12237) := x"0020";
    tmp(12238) := x"0020";
    tmp(12239) := x"0020";
    tmp(12240) := x"0000";
    tmp(12241) := x"0041";
    tmp(12242) := x"0041";
    tmp(12243) := x"0041";
    tmp(12244) := x"0061";
    tmp(12245) := x"0061";
    tmp(12246) := x"0041";
    tmp(12247) := x"0061";
    tmp(12248) := x"0861";
    tmp(12249) := x"0861";
    tmp(12250) := x"0861";
    tmp(12251) := x"10a1";
    tmp(12252) := x"20e0";
    tmp(12253) := x"3120";
    tmp(12254) := x"4960";
    tmp(12255) := x"59a0";
    tmp(12256) := x"61a0";
    tmp(12257) := x"6a00";
    tmp(12258) := x"7200";
    tmp(12259) := x"7200";
    tmp(12260) := x"7200";
    tmp(12261) := x"71e0";
    tmp(12262) := x"71e0";
    tmp(12263) := x"71e0";
    tmp(12264) := x"71c0";
    tmp(12265) := x"71e0";
    tmp(12266) := x"71e0";
    tmp(12267) := x"79e0";
    tmp(12268) := x"71e0";
    tmp(12269) := x"79e0";
    tmp(12270) := x"7a00";
    tmp(12271) := x"8a40";
    tmp(12272) := x"8a40";
    tmp(12273) := x"8a60";
    tmp(12274) := x"8a60";
    tmp(12275) := x"8240";
    tmp(12276) := x"8a60";
    tmp(12277) := x"7a40";
    tmp(12278) := x"6a40";
    tmp(12279) := x"6221";
    tmp(12280) := x"7281";
    tmp(12281) := x"7aa1";
    tmp(12282) := x"82a1";
    tmp(12283) := x"7aa2";
    tmp(12284) := x"8ac1";
    tmp(12285) := x"9ac0";
    tmp(12286) := x"8aa0";
    tmp(12287) := x"59e0";
    tmp(12288) := x"28e0";
    tmp(12289) := x"0820";
    tmp(12290) := x"0820";
    tmp(12291) := x"0820";
    tmp(12292) := x"0820";
    tmp(12293) := x"0820";
    tmp(12294) := x"0820";
    tmp(12295) := x"0820";
    tmp(12296) := x"0820";
    tmp(12297) := x"0820";
    tmp(12298) := x"0820";
    tmp(12299) := x"0820";
    tmp(12300) := x"0820";
    tmp(12301) := x"0820";
    tmp(12302) := x"0820";
    tmp(12303) := x"0820";
    tmp(12304) := x"0820";
    tmp(12305) := x"0820";
    tmp(12306) := x"0820";
    tmp(12307) := x"0820";
    tmp(12308) := x"0820";
    tmp(12309) := x"0840";
    tmp(12310) := x"0820";
    tmp(12311) := x"0820";
    tmp(12312) := x"0820";
    tmp(12313) := x"0820";
    tmp(12314) := x"0820";
    tmp(12315) := x"0820";
    tmp(12316) := x"0820";
    tmp(12317) := x"0840";
    tmp(12318) := x"0860";
    tmp(12319) := x"0840";
    tmp(12320) := x"0020";
    tmp(12321) := x"0020";
    tmp(12322) := x"0020";
    tmp(12323) := x"0020";
    tmp(12324) := x"0000";
    tmp(12325) := x"0000";
    tmp(12326) := x"0000";
    tmp(12327) := x"0000";
    tmp(12328) := x"0000";
    tmp(12329) := x"0000";
    tmp(12330) := x"0000";
    tmp(12331) := x"0000";
    tmp(12332) := x"0000";
    tmp(12333) := x"0000";
    tmp(12334) := x"0000";
    tmp(12335) := x"0000";
    tmp(12336) := x"0000";
    tmp(12337) := x"0000";
    tmp(12338) := x"18a2";
    tmp(12339) := x"1082";
    tmp(12340) := x"0000";
    tmp(12341) := x"0000";
    tmp(12342) := x"0000";
    tmp(12343) := x"0000";
    tmp(12344) := x"0000";
    tmp(12345) := x"0000";
    tmp(12346) := x"0000";
    tmp(12347) := x"0000";
    tmp(12348) := x"0000";
    tmp(12349) := x"0000";
    tmp(12350) := x"0000";
    tmp(12351) := x"0000";
    tmp(12352) := x"0000";
    tmp(12353) := x"0000";
    tmp(12354) := x"0000";
    tmp(12355) := x"0000";
    tmp(12356) := x"0000";
    tmp(12357) := x"0000";
    tmp(12358) := x"0000";
    tmp(12359) := x"0000";
    tmp(12360) := x"0000";
    tmp(12361) := x"1082";
    tmp(12362) := x"6b0c";
    tmp(12363) := x"5a29";
    tmp(12364) := x"3925";
    tmp(12365) := x"abf0";
    tmp(12366) := x"9bb0";
    tmp(12367) := x"93af";
    tmp(12368) := x"9bd0";
    tmp(12369) := x"9baf";
    tmp(12370) := x"9bcf";
    tmp(12371) := x"9c11";
    tmp(12372) := x"a412";
    tmp(12373) := x"ac72";
    tmp(12374) := x"ac72";
    tmp(12375) := x"b473";
    tmp(12376) := x"ac12";
    tmp(12377) := x"830e";
    tmp(12378) := x"6a4b";
    tmp(12379) := x"82cd";
    tmp(12380) := x"8b0d";
    tmp(12381) := x"934d";
    tmp(12382) := x"6a4a";
    tmp(12383) := x"4986";
    tmp(12384) := x"3925";
    tmp(12385) := x"20a3";
    tmp(12386) := x"2082";
    tmp(12387) := x"38e4";
    tmp(12388) := x"bbaf";
    tmp(12389) := x"e536";
    tmp(12390) := x"e512";
    tmp(12391) := x"9bcc";
    tmp(12392) := x"0020";
    tmp(12393) := x"0860";
    tmp(12394) := x"0880";
    tmp(12395) := x"0840";
    tmp(12396) := x"10e0";
    tmp(12397) := x"10e0";
    tmp(12398) := x"0860";
    tmp(12399) := x"0860";
    tmp(12400) := x"0860";
    tmp(12401) := x"0860";
    tmp(12402) := x"0860";
    tmp(12403) := x"0040";
    tmp(12404) := x"0040";
    tmp(12405) := x"0040";
    tmp(12406) := x"0040";
    tmp(12407) := x"0040";
    tmp(12408) := x"0040";
    tmp(12409) := x"0040";
    tmp(12410) := x"0040";
    tmp(12411) := x"0040";
    tmp(12412) := x"0060";
    tmp(12413) := x"0060";
    tmp(12414) := x"0060";
    tmp(12415) := x"0060";
    tmp(12416) := x"0860";
    tmp(12417) := x"0860";
    tmp(12418) := x"0880";
    tmp(12419) := x"0880";
    tmp(12420) := x"0880";
    tmp(12421) := x"08a0";
    tmp(12422) := x"08a0";
    tmp(12423) := x"08a0";
    tmp(12424) := x"08a0";
    tmp(12425) := x"08a0";
    tmp(12426) := x"08a0";
    tmp(12427) := x"08a0";
    tmp(12428) := x"08a0";
    tmp(12429) := x"08a0";
    tmp(12430) := x"08a0";
    tmp(12431) := x"00a0";
    tmp(12432) := x"08a0";
    tmp(12433) := x"0080";
    tmp(12434) := x"0080";
    tmp(12435) := x"0080";
    tmp(12436) := x"0060";
    tmp(12437) := x"0000";
    tmp(12438) := x"0000";
    tmp(12439) := x"0000";
    tmp(12440) := x"0000";
    tmp(12441) := x"0000";
    tmp(12442) := x"0000";
    tmp(12443) := x"0000";
    tmp(12444) := x"0000";
    tmp(12445) := x"0000";
    tmp(12446) := x"0000";
    tmp(12447) := x"0000";
    tmp(12448) := x"0000";
    tmp(12449) := x"0000";
    tmp(12450) := x"0000";
    tmp(12451) := x"0000";
    tmp(12452) := x"0000";
    tmp(12453) := x"0000";
    tmp(12454) := x"0000";
    tmp(12455) := x"0000";
    tmp(12456) := x"0000";
    tmp(12457) := x"0000";
    tmp(12458) := x"0000";
    tmp(12459) := x"0000";
    tmp(12460) := x"0000";
    tmp(12461) := x"0000";
    tmp(12462) := x"0000";
    tmp(12463) := x"0000";
    tmp(12464) := x"0000";
    tmp(12465) := x"0000";
    tmp(12466) := x"0000";
    tmp(12467) := x"0000";
    tmp(12468) := x"0000";
    tmp(12469) := x"0000";
    tmp(12470) := x"0000";
    tmp(12471) := x"0000";
    tmp(12472) := x"0000";
    tmp(12473) := x"0000";
    tmp(12474) := x"0000";
    tmp(12475) := x"0000";
    tmp(12476) := x"0000";
    tmp(12477) := x"0020";
    tmp(12478) := x"0020";
    tmp(12479) := x"0020";
    tmp(12480) := x"0000";
    tmp(12481) := x"0041";
    tmp(12482) := x"0041";
    tmp(12483) := x"0041";
    tmp(12484) := x"0041";
    tmp(12485) := x"0041";
    tmp(12486) := x"0041";
    tmp(12487) := x"0041";
    tmp(12488) := x"0041";
    tmp(12489) := x"0861";
    tmp(12490) := x"0861";
    tmp(12491) := x"0840";
    tmp(12492) := x"1060";
    tmp(12493) := x"28c0";
    tmp(12494) := x"4140";
    tmp(12495) := x"5180";
    tmp(12496) := x"69e0";
    tmp(12497) := x"7200";
    tmp(12498) := x"7200";
    tmp(12499) := x"7a20";
    tmp(12500) := x"8200";
    tmp(12501) := x"8200";
    tmp(12502) := x"8a20";
    tmp(12503) := x"8a00";
    tmp(12504) := x"81e0";
    tmp(12505) := x"81e0";
    tmp(12506) := x"8200";
    tmp(12507) := x"8200";
    tmp(12508) := x"9240";
    tmp(12509) := x"9a60";
    tmp(12510) := x"9a80";
    tmp(12511) := x"9280";
    tmp(12512) := x"9aa0";
    tmp(12513) := x"a2c0";
    tmp(12514) := x"9aa0";
    tmp(12515) := x"9aa0";
    tmp(12516) := x"9aa0";
    tmp(12517) := x"9aa0";
    tmp(12518) := x"9ac0";
    tmp(12519) := x"9ac0";
    tmp(12520) := x"a300";
    tmp(12521) := x"ab00";
    tmp(12522) := x"ab00";
    tmp(12523) := x"b340";
    tmp(12524) := x"bb20";
    tmp(12525) := x"b320";
    tmp(12526) := x"b340";
    tmp(12527) := x"b300";
    tmp(12528) := x"8260";
    tmp(12529) := x"3920";
    tmp(12530) := x"28e0";
    tmp(12531) := x"20c0";
    tmp(12532) := x"1880";
    tmp(12533) := x"0840";
    tmp(12534) := x"0820";
    tmp(12535) := x"0820";
    tmp(12536) := x"0820";
    tmp(12537) := x"0820";
    tmp(12538) := x"0820";
    tmp(12539) := x"0820";
    tmp(12540) := x"0820";
    tmp(12541) := x"0820";
    tmp(12542) := x"0820";
    tmp(12543) := x"0820";
    tmp(12544) := x"0820";
    tmp(12545) := x"0820";
    tmp(12546) := x"0820";
    tmp(12547) := x"0820";
    tmp(12548) := x"0820";
    tmp(12549) := x"0820";
    tmp(12550) := x"0820";
    tmp(12551) := x"0820";
    tmp(12552) := x"0820";
    tmp(12553) := x"0840";
    tmp(12554) := x"0860";
    tmp(12555) := x"10a0";
    tmp(12556) := x"1081";
    tmp(12557) := x"0840";
    tmp(12558) := x"0820";
    tmp(12559) := x"0020";
    tmp(12560) := x"0000";
    tmp(12561) := x"0000";
    tmp(12562) := x"0000";
    tmp(12563) := x"0000";
    tmp(12564) := x"0000";
    tmp(12565) := x"0000";
    tmp(12566) := x"0000";
    tmp(12567) := x"0000";
    tmp(12568) := x"0000";
    tmp(12569) := x"0000";
    tmp(12570) := x"0000";
    tmp(12571) := x"0000";
    tmp(12572) := x"0000";
    tmp(12573) := x"0000";
    tmp(12574) := x"0000";
    tmp(12575) := x"0000";
    tmp(12576) := x"0000";
    tmp(12577) := x"0000";
    tmp(12578) := x"0841";
    tmp(12579) := x"3165";
    tmp(12580) := x"1082";
    tmp(12581) := x"0000";
    tmp(12582) := x"0000";
    tmp(12583) := x"0000";
    tmp(12584) := x"0000";
    tmp(12585) := x"0000";
    tmp(12586) := x"0000";
    tmp(12587) := x"0000";
    tmp(12588) := x"0000";
    tmp(12589) := x"0000";
    tmp(12590) := x"0000";
    tmp(12591) := x"0000";
    tmp(12592) := x"0000";
    tmp(12593) := x"0000";
    tmp(12594) := x"0000";
    tmp(12595) := x"0000";
    tmp(12596) := x"0000";
    tmp(12597) := x"0000";
    tmp(12598) := x"0000";
    tmp(12599) := x"0820";
    tmp(12600) := x"2924";
    tmp(12601) := x"7b6e";
    tmp(12602) := x"c578";
    tmp(12603) := x"8b70";
    tmp(12604) := x"4145";
    tmp(12605) := x"930d";
    tmp(12606) := x"ccf6";
    tmp(12607) := x"bc95";
    tmp(12608) := x"bc74";
    tmp(12609) := x"9b70";
    tmp(12610) := x"b3f2";
    tmp(12611) := x"bc74";
    tmp(12612) := x"bcb6";
    tmp(12613) := x"b453";
    tmp(12614) := x"ac12";
    tmp(12615) := x"93b2";
    tmp(12616) := x"9391";
    tmp(12617) := x"6a6b";
    tmp(12618) := x"726b";
    tmp(12619) := x"8b2e";
    tmp(12620) := x"b431";
    tmp(12621) := x"4165";
    tmp(12622) := x"0821";
    tmp(12623) := x"0820";
    tmp(12624) := x"0841";
    tmp(12625) := x"0841";
    tmp(12626) := x"0800";
    tmp(12627) := x"28a2";
    tmp(12628) := x"cc71";
    tmp(12629) := x"e491";
    tmp(12630) := x"fef8";
    tmp(12631) := x"20c2";
    tmp(12632) := x"0020";
    tmp(12633) := x"0860";
    tmp(12634) := x"10c0";
    tmp(12635) := x"10c0";
    tmp(12636) := x"1940";
    tmp(12637) := x"1120";
    tmp(12638) := x"0880";
    tmp(12639) := x"0060";
    tmp(12640) := x"0860";
    tmp(12641) := x"0060";
    tmp(12642) := x"0040";
    tmp(12643) := x"0040";
    tmp(12644) := x"0040";
    tmp(12645) := x"0040";
    tmp(12646) := x"0040";
    tmp(12647) := x"0040";
    tmp(12648) := x"0040";
    tmp(12649) := x"0040";
    tmp(12650) := x"0040";
    tmp(12651) := x"0040";
    tmp(12652) := x"0040";
    tmp(12653) := x"0040";
    tmp(12654) := x"0040";
    tmp(12655) := x"0840";
    tmp(12656) := x"0860";
    tmp(12657) := x"0860";
    tmp(12658) := x"0860";
    tmp(12659) := x"0860";
    tmp(12660) := x"0860";
    tmp(12661) := x"0880";
    tmp(12662) := x"0880";
    tmp(12663) := x"0880";
    tmp(12664) := x"0880";
    tmp(12665) := x"08a0";
    tmp(12666) := x"08a0";
    tmp(12667) := x"08a0";
    tmp(12668) := x"08a0";
    tmp(12669) := x"0880";
    tmp(12670) := x"0880";
    tmp(12671) := x"0080";
    tmp(12672) := x"0080";
    tmp(12673) := x"0080";
    tmp(12674) := x"0080";
    tmp(12675) := x"0080";
    tmp(12676) := x"0080";
    tmp(12677) := x"0000";
    tmp(12678) := x"0000";
    tmp(12679) := x"0000";
    tmp(12680) := x"0000";
    tmp(12681) := x"0000";
    tmp(12682) := x"0000";
    tmp(12683) := x"0000";
    tmp(12684) := x"0000";
    tmp(12685) := x"0000";
    tmp(12686) := x"0000";
    tmp(12687) := x"0000";
    tmp(12688) := x"0000";
    tmp(12689) := x"0000";
    tmp(12690) := x"0000";
    tmp(12691) := x"0000";
    tmp(12692) := x"0000";
    tmp(12693) := x"0000";
    tmp(12694) := x"0000";
    tmp(12695) := x"0000";
    tmp(12696) := x"0000";
    tmp(12697) := x"0000";
    tmp(12698) := x"0000";
    tmp(12699) := x"0000";
    tmp(12700) := x"0000";
    tmp(12701) := x"0000";
    tmp(12702) := x"0000";
    tmp(12703) := x"0000";
    tmp(12704) := x"0000";
    tmp(12705) := x"0000";
    tmp(12706) := x"0000";
    tmp(12707) := x"0000";
    tmp(12708) := x"0000";
    tmp(12709) := x"0000";
    tmp(12710) := x"0000";
    tmp(12711) := x"0000";
    tmp(12712) := x"0000";
    tmp(12713) := x"0000";
    tmp(12714) := x"0000";
    tmp(12715) := x"0000";
    tmp(12716) := x"0000";
    tmp(12717) := x"0020";
    tmp(12718) := x"0020";
    tmp(12719) := x"0020";
    tmp(12720) := x"0000";
    tmp(12721) := x"0020";
    tmp(12722) := x"0020";
    tmp(12723) := x"0020";
    tmp(12724) := x"0020";
    tmp(12725) := x"0020";
    tmp(12726) := x"0041";
    tmp(12727) := x"0861";
    tmp(12728) := x"1080";
    tmp(12729) := x"18a0";
    tmp(12730) := x"20c0";
    tmp(12731) := x"2900";
    tmp(12732) := x"3100";
    tmp(12733) := x"30e0";
    tmp(12734) := x"3900";
    tmp(12735) := x"59a0";
    tmp(12736) := x"69e0";
    tmp(12737) := x"8220";
    tmp(12738) := x"8240";
    tmp(12739) := x"8a20";
    tmp(12740) := x"9240";
    tmp(12741) := x"9260";
    tmp(12742) := x"9260";
    tmp(12743) := x"9240";
    tmp(12744) := x"9220";
    tmp(12745) := x"9200";
    tmp(12746) := x"9220";
    tmp(12747) := x"9240";
    tmp(12748) := x"9a60";
    tmp(12749) := x"9a80";
    tmp(12750) := x"a2a0";
    tmp(12751) := x"a2a0";
    tmp(12752) := x"a2a0";
    tmp(12753) := x"9a80";
    tmp(12754) := x"aaa0";
    tmp(12755) := x"a2a0";
    tmp(12756) := x"a2a0";
    tmp(12757) := x"aac0";
    tmp(12758) := x"aac0";
    tmp(12759) := x"b300";
    tmp(12760) := x"bb40";
    tmp(12761) := x"b340";
    tmp(12762) := x"bb40";
    tmp(12763) := x"bb40";
    tmp(12764) := x"c380";
    tmp(12765) := x"c340";
    tmp(12766) := x"c340";
    tmp(12767) := x"bb40";
    tmp(12768) := x"bb40";
    tmp(12769) := x"b320";
    tmp(12770) := x"ab00";
    tmp(12771) := x"a2c0";
    tmp(12772) := x"9aa0";
    tmp(12773) := x"7a60";
    tmp(12774) := x"4140";
    tmp(12775) := x"1880";
    tmp(12776) := x"0840";
    tmp(12777) := x"0820";
    tmp(12778) := x"0820";
    tmp(12779) := x"0820";
    tmp(12780) := x"0820";
    tmp(12781) := x"0820";
    tmp(12782) := x"0820";
    tmp(12783) := x"0820";
    tmp(12784) := x"0820";
    tmp(12785) := x"0820";
    tmp(12786) := x"0820";
    tmp(12787) := x"1060";
    tmp(12788) := x"20c0";
    tmp(12789) := x"3920";
    tmp(12790) := x"51a0";
    tmp(12791) := x"5a01";
    tmp(12792) := x"49c1";
    tmp(12793) := x"2961";
    tmp(12794) := x"2120";
    tmp(12795) := x"18e0";
    tmp(12796) := x"0860";
    tmp(12797) := x"0020";
    tmp(12798) := x"0000";
    tmp(12799) := x"0000";
    tmp(12800) := x"0000";
    tmp(12801) := x"0000";
    tmp(12802) := x"0000";
    tmp(12803) := x"0000";
    tmp(12804) := x"0000";
    tmp(12805) := x"0000";
    tmp(12806) := x"0000";
    tmp(12807) := x"0000";
    tmp(12808) := x"0000";
    tmp(12809) := x"0000";
    tmp(12810) := x"0000";
    tmp(12811) := x"0000";
    tmp(12812) := x"0000";
    tmp(12813) := x"0000";
    tmp(12814) := x"0000";
    tmp(12815) := x"0000";
    tmp(12816) := x"0000";
    tmp(12817) := x"0000";
    tmp(12818) := x"0840";
    tmp(12819) := x"20e3";
    tmp(12820) := x"2904";
    tmp(12821) := x"2124";
    tmp(12822) := x"1061";
    tmp(12823) := x"0000";
    tmp(12824) := x"0000";
    tmp(12825) := x"0000";
    tmp(12826) := x"0000";
    tmp(12827) := x"0000";
    tmp(12828) := x"0000";
    tmp(12829) := x"0000";
    tmp(12830) := x"0000";
    tmp(12831) := x"0000";
    tmp(12832) := x"0000";
    tmp(12833) := x"0000";
    tmp(12834) := x"0000";
    tmp(12835) := x"0000";
    tmp(12836) := x"0020";
    tmp(12837) := x"1082";
    tmp(12838) := x"3145";
    tmp(12839) := x"732d";
    tmp(12840) := x"8b8f";
    tmp(12841) := x"bcf5";
    tmp(12842) := x"bcf7";
    tmp(12843) := x"a3f2";
    tmp(12844) := x"4945";
    tmp(12845) := x"8a8b";
    tmp(12846) := x"d4f6";
    tmp(12847) := x"dd9a";
    tmp(12848) := x"a3d2";
    tmp(12849) := x"9390";
    tmp(12850) := x"6a2a";
    tmp(12851) := x"82ad";
    tmp(12852) := x"728c";
    tmp(12853) := x"8b2f";
    tmp(12854) := x"a3d2";
    tmp(12855) := x"6a4b";
    tmp(12856) := x"6a4a";
    tmp(12857) := x"8b0d";
    tmp(12858) := x"7aac";
    tmp(12859) := x"8b0d";
    tmp(12860) := x"9b6f";
    tmp(12861) := x"5a08";
    tmp(12862) := x"0841";
    tmp(12863) := x"0000";
    tmp(12864) := x"0000";
    tmp(12865) := x"0820";
    tmp(12866) := x"1861";
    tmp(12867) := x"59a6";
    tmp(12868) := x"cc72";
    tmp(12869) := x"fd33";
    tmp(12870) := x"c48f";
    tmp(12871) := x"0820";
    tmp(12872) := x"0840";
    tmp(12873) := x"0880";
    tmp(12874) := x"10e0";
    tmp(12875) := x"1900";
    tmp(12876) := x"2160";
    tmp(12877) := x"21c0";
    tmp(12878) := x"08a0";
    tmp(12879) := x"0060";
    tmp(12880) := x"0860";
    tmp(12881) := x"0860";
    tmp(12882) := x"0040";
    tmp(12883) := x"0040";
    tmp(12884) := x"0040";
    tmp(12885) := x"0040";
    tmp(12886) := x"0040";
    tmp(12887) := x"0040";
    tmp(12888) := x"0040";
    tmp(12889) := x"0040";
    tmp(12890) := x"0040";
    tmp(12891) := x"0040";
    tmp(12892) := x"0040";
    tmp(12893) := x"0040";
    tmp(12894) := x"0840";
    tmp(12895) := x"0840";
    tmp(12896) := x"0840";
    tmp(12897) := x"0840";
    tmp(12898) := x"0860";
    tmp(12899) := x"0860";
    tmp(12900) := x"0860";
    tmp(12901) := x"0860";
    tmp(12902) := x"0860";
    tmp(12903) := x"0860";
    tmp(12904) := x"0860";
    tmp(12905) := x"0880";
    tmp(12906) := x"0880";
    tmp(12907) := x"0880";
    tmp(12908) := x"0880";
    tmp(12909) := x"0880";
    tmp(12910) := x"0880";
    tmp(12911) := x"0080";
    tmp(12912) := x"0880";
    tmp(12913) := x"0080";
    tmp(12914) := x"0080";
    tmp(12915) := x"0080";
    tmp(12916) := x"0080";
    tmp(12917) := x"0000";
    tmp(12918) := x"0000";
    tmp(12919) := x"0000";
    tmp(12920) := x"0000";
    tmp(12921) := x"0000";
    tmp(12922) := x"0000";
    tmp(12923) := x"0000";
    tmp(12924) := x"0000";
    tmp(12925) := x"0000";
    tmp(12926) := x"0000";
    tmp(12927) := x"0000";
    tmp(12928) := x"0000";
    tmp(12929) := x"0000";
    tmp(12930) := x"0000";
    tmp(12931) := x"0000";
    tmp(12932) := x"0000";
    tmp(12933) := x"0000";
    tmp(12934) := x"0000";
    tmp(12935) := x"0000";
    tmp(12936) := x"0000";
    tmp(12937) := x"0000";
    tmp(12938) := x"0000";
    tmp(12939) := x"0000";
    tmp(12940) := x"0000";
    tmp(12941) := x"0000";
    tmp(12942) := x"0000";
    tmp(12943) := x"0000";
    tmp(12944) := x"0000";
    tmp(12945) := x"0000";
    tmp(12946) := x"0000";
    tmp(12947) := x"0000";
    tmp(12948) := x"0000";
    tmp(12949) := x"0000";
    tmp(12950) := x"0000";
    tmp(12951) := x"0000";
    tmp(12952) := x"0000";
    tmp(12953) := x"0000";
    tmp(12954) := x"0000";
    tmp(12955) := x"0000";
    tmp(12956) := x"0000";
    tmp(12957) := x"0000";
    tmp(12958) := x"0020";
    tmp(12959) := x"0020";
    tmp(12960) := x"0000";
    tmp(12961) := x"0020";
    tmp(12962) := x"0020";
    tmp(12963) := x"0020";
    tmp(12964) := x"0020";
    tmp(12965) := x"0020";
    tmp(12966) := x"0880";
    tmp(12967) := x"20e0";
    tmp(12968) := x"3120";
    tmp(12969) := x"3940";
    tmp(12970) := x"4960";
    tmp(12971) := x"51a0";
    tmp(12972) := x"6a00";
    tmp(12973) := x"7220";
    tmp(12974) := x"7a40";
    tmp(12975) := x"7a20";
    tmp(12976) := x"7a20";
    tmp(12977) := x"8a40";
    tmp(12978) := x"9260";
    tmp(12979) := x"9a60";
    tmp(12980) := x"9a60";
    tmp(12981) := x"9a60";
    tmp(12982) := x"9a60";
    tmp(12983) := x"9a40";
    tmp(12984) := x"9a40";
    tmp(12985) := x"9a40";
    tmp(12986) := x"9a60";
    tmp(12987) := x"a280";
    tmp(12988) := x"a280";
    tmp(12989) := x"9a80";
    tmp(12990) := x"9a80";
    tmp(12991) := x"a280";
    tmp(12992) := x"9a80";
    tmp(12993) := x"a2a0";
    tmp(12994) := x"a2a0";
    tmp(12995) := x"aaa0";
    tmp(12996) := x"aac0";
    tmp(12997) := x"aac0";
    tmp(12998) := x"aac0";
    tmp(12999) := x"b320";
    tmp(13000) := x"bb40";
    tmp(13001) := x"bb20";
    tmp(13002) := x"c340";
    tmp(13003) := x"c360";
    tmp(13004) := x"c360";
    tmp(13005) := x"d380";
    tmp(13006) := x"cb60";
    tmp(13007) := x"cb40";
    tmp(13008) := x"bb00";
    tmp(13009) := x"db80";
    tmp(13010) := x"d340";
    tmp(13011) := x"cb40";
    tmp(13012) := x"cb40";
    tmp(13013) := x"cb40";
    tmp(13014) := x"c340";
    tmp(13015) := x"ab00";
    tmp(13016) := x"8260";
    tmp(13017) := x"4980";
    tmp(13018) := x"28c0";
    tmp(13019) := x"20a0";
    tmp(13020) := x"20a0";
    tmp(13021) := x"1880";
    tmp(13022) := x"1860";
    tmp(13023) := x"1060";
    tmp(13024) := x"1060";
    tmp(13025) := x"20a0";
    tmp(13026) := x"5180";
    tmp(13027) := x"8a80";
    tmp(13028) := x"a2c0";
    tmp(13029) := x"aac0";
    tmp(13030) := x"aac0";
    tmp(13031) := x"7a20";
    tmp(13032) := x"51a0";
    tmp(13033) := x"3140";
    tmp(13034) := x"18e0";
    tmp(13035) := x"1060";
    tmp(13036) := x"0820";
    tmp(13037) := x"0020";
    tmp(13038) := x"0000";
    tmp(13039) := x"0000";
    tmp(13040) := x"0000";
    tmp(13041) := x"0000";
    tmp(13042) := x"0000";
    tmp(13043) := x"0000";
    tmp(13044) := x"0000";
    tmp(13045) := x"0000";
    tmp(13046) := x"0000";
    tmp(13047) := x"0000";
    tmp(13048) := x"0000";
    tmp(13049) := x"0000";
    tmp(13050) := x"0000";
    tmp(13051) := x"0000";
    tmp(13052) := x"0000";
    tmp(13053) := x"0000";
    tmp(13054) := x"0000";
    tmp(13055) := x"0000";
    tmp(13056) := x"0000";
    tmp(13057) := x"0000";
    tmp(13058) := x"0820";
    tmp(13059) := x"2904";
    tmp(13060) := x"2104";
    tmp(13061) := x"2105";
    tmp(13062) := x"2945";
    tmp(13063) := x"31a6";
    tmp(13064) := x"2924";
    tmp(13065) := x"10a2";
    tmp(13066) := x"1082";
    tmp(13067) := x"10a2";
    tmp(13068) := x"10a2";
    tmp(13069) := x"18c3";
    tmp(13070) := x"20e4";
    tmp(13071) := x"2104";
    tmp(13072) := x"3165";
    tmp(13073) := x"39c7";
    tmp(13074) := x"41e8";
    tmp(13075) := x"5acb";
    tmp(13076) := x"734e";
    tmp(13077) := x"732d";
    tmp(13078) := x"a452";
    tmp(13079) := x"bcb6";
    tmp(13080) := x"9bb1";
    tmp(13081) := x"ac54";
    tmp(13082) := x"c4f8";
    tmp(13083) := x"b413";
    tmp(13084) := x"7229";
    tmp(13085) := x"8aab";
    tmp(13086) := x"930e";
    tmp(13087) := x"c4b6";
    tmp(13088) := x"ac55";
    tmp(13089) := x"8b50";
    tmp(13090) := x"934f";
    tmp(13091) := x"49a7";
    tmp(13092) := x"8b0d";
    tmp(13093) := x"9bb1";
    tmp(13094) := x"49a8";
    tmp(13095) := x"6a6b";
    tmp(13096) := x"8b2e";
    tmp(13097) := x"82ac";
    tmp(13098) := x"6a0a";
    tmp(13099) := x"82ed";
    tmp(13100) := x"934f";
    tmp(13101) := x"bc72";
    tmp(13102) := x"6a69";
    tmp(13103) := x"51a6";
    tmp(13104) := x"49a6";
    tmp(13105) := x"4164";
    tmp(13106) := x"7a89";
    tmp(13107) := x"cc51";
    tmp(13108) := x"cc50";
    tmp(13109) := x"fed7";
    tmp(13110) := x"28c2";
    tmp(13111) := x"0840";
    tmp(13112) := x"0860";
    tmp(13113) := x"08a0";
    tmp(13114) := x"10e0";
    tmp(13115) := x"1920";
    tmp(13116) := x"29a0";
    tmp(13117) := x"2a00";
    tmp(13118) := x"08c0";
    tmp(13119) := x"0860";
    tmp(13120) := x"0860";
    tmp(13121) := x"0860";
    tmp(13122) := x"0060";
    tmp(13123) := x"0860";
    tmp(13124) := x"0040";
    tmp(13125) := x"0040";
    tmp(13126) := x"0040";
    tmp(13127) := x"0040";
    tmp(13128) := x"0040";
    tmp(13129) := x"0040";
    tmp(13130) := x"0040";
    tmp(13131) := x"0040";
    tmp(13132) := x"0040";
    tmp(13133) := x"0040";
    tmp(13134) := x"0840";
    tmp(13135) := x"0840";
    tmp(13136) := x"0840";
    tmp(13137) := x"0840";
    tmp(13138) := x"0840";
    tmp(13139) := x"0840";
    tmp(13140) := x"0840";
    tmp(13141) := x"0860";
    tmp(13142) := x"0860";
    tmp(13143) := x"0860";
    tmp(13144) := x"0860";
    tmp(13145) := x"0860";
    tmp(13146) := x"0860";
    tmp(13147) := x"0860";
    tmp(13148) := x"0860";
    tmp(13149) := x"0880";
    tmp(13150) := x"0880";
    tmp(13151) := x"0880";
    tmp(13152) := x"0080";
    tmp(13153) := x"0080";
    tmp(13154) := x"0060";
    tmp(13155) := x"0080";
    tmp(13156) := x"0080";
    tmp(13157) := x"0000";
    tmp(13158) := x"0000";
    tmp(13159) := x"0000";
    tmp(13160) := x"0000";
    tmp(13161) := x"0000";
    tmp(13162) := x"0000";
    tmp(13163) := x"0000";
    tmp(13164) := x"0000";
    tmp(13165) := x"0000";
    tmp(13166) := x"0000";
    tmp(13167) := x"0000";
    tmp(13168) := x"0000";
    tmp(13169) := x"0000";
    tmp(13170) := x"0000";
    tmp(13171) := x"0000";
    tmp(13172) := x"0000";
    tmp(13173) := x"0000";
    tmp(13174) := x"0000";
    tmp(13175) := x"0000";
    tmp(13176) := x"0000";
    tmp(13177) := x"0000";
    tmp(13178) := x"0000";
    tmp(13179) := x"0000";
    tmp(13180) := x"0000";
    tmp(13181) := x"0000";
    tmp(13182) := x"0000";
    tmp(13183) := x"0000";
    tmp(13184) := x"0000";
    tmp(13185) := x"0000";
    tmp(13186) := x"0000";
    tmp(13187) := x"0000";
    tmp(13188) := x"0000";
    tmp(13189) := x"0000";
    tmp(13190) := x"0000";
    tmp(13191) := x"0000";
    tmp(13192) := x"0000";
    tmp(13193) := x"0000";
    tmp(13194) := x"0000";
    tmp(13195) := x"0000";
    tmp(13196) := x"0000";
    tmp(13197) := x"0000";
    tmp(13198) := x"0020";
    tmp(13199) := x"0020";
    tmp(13200) := x"0820";
    tmp(13201) := x"49c0";
    tmp(13202) := x"3940";
    tmp(13203) := x"28e0";
    tmp(13204) := x"18a0";
    tmp(13205) := x"20c0";
    tmp(13206) := x"3960";
    tmp(13207) := x"59c0";
    tmp(13208) := x"7220";
    tmp(13209) := x"8260";
    tmp(13210) := x"8260";
    tmp(13211) := x"8a60";
    tmp(13212) := x"9280";
    tmp(13213) := x"8a60";
    tmp(13214) := x"9280";
    tmp(13215) := x"9a80";
    tmp(13216) := x"a280";
    tmp(13217) := x"a280";
    tmp(13218) := x"aac0";
    tmp(13219) := x"aaa0";
    tmp(13220) := x"a260";
    tmp(13221) := x"a260";
    tmp(13222) := x"a280";
    tmp(13223) := x"aa80";
    tmp(13224) := x"a280";
    tmp(13225) := x"a260";
    tmp(13226) := x"a260";
    tmp(13227) := x"a280";
    tmp(13228) := x"a280";
    tmp(13229) := x"a280";
    tmp(13230) := x"a280";
    tmp(13231) := x"a280";
    tmp(13232) := x"a280";
    tmp(13233) := x"aaa0";
    tmp(13234) := x"aaa0";
    tmp(13235) := x"aac0";
    tmp(13236) := x"aac0";
    tmp(13237) := x"aac0";
    tmp(13238) := x"aac0";
    tmp(13239) := x"b2e0";
    tmp(13240) := x"b2e0";
    tmp(13241) := x"bb00";
    tmp(13242) := x"bb00";
    tmp(13243) := x"c340";
    tmp(13244) := x"c340";
    tmp(13245) := x"cb40";
    tmp(13246) := x"bb00";
    tmp(13247) := x"c2e0";
    tmp(13248) := x"bac0";
    tmp(13249) := x"bac0";
    tmp(13250) := x"bac0";
    tmp(13251) := x"bae0";
    tmp(13252) := x"bb00";
    tmp(13253) := x"c300";
    tmp(13254) := x"c300";
    tmp(13255) := x"c320";
    tmp(13256) := x"c320";
    tmp(13257) := x"bb00";
    tmp(13258) := x"c340";
    tmp(13259) := x"b320";
    tmp(13260) := x"b340";
    tmp(13261) := x"b340";
    tmp(13262) := x"b320";
    tmp(13263) := x"b360";
    tmp(13264) := x"b360";
    tmp(13265) := x"bb80";
    tmp(13266) := x"ab00";
    tmp(13267) := x"9a80";
    tmp(13268) := x"9a60";
    tmp(13269) := x"9a60";
    tmp(13270) := x"9260";
    tmp(13271) := x"79e0";
    tmp(13272) := x"4960";
    tmp(13273) := x"3120";
    tmp(13274) := x"18a0";
    tmp(13275) := x"0840";
    tmp(13276) := x"0020";
    tmp(13277) := x"0000";
    tmp(13278) := x"0020";
    tmp(13279) := x"0000";
    tmp(13280) := x"0000";
    tmp(13281) := x"0000";
    tmp(13282) := x"0000";
    tmp(13283) := x"0000";
    tmp(13284) := x"0000";
    tmp(13285) := x"0000";
    tmp(13286) := x"0000";
    tmp(13287) := x"0000";
    tmp(13288) := x"0000";
    tmp(13289) := x"0000";
    tmp(13290) := x"0000";
    tmp(13291) := x"0000";
    tmp(13292) := x"0000";
    tmp(13293) := x"0000";
    tmp(13294) := x"0000";
    tmp(13295) := x"0000";
    tmp(13296) := x"0000";
    tmp(13297) := x"0000";
    tmp(13298) := x"0820";
    tmp(13299) := x"28e4";
    tmp(13300) := x"3987";
    tmp(13301) := x"2926";
    tmp(13302) := x"2926";
    tmp(13303) := x"3146";
    tmp(13304) := x"3187";
    tmp(13305) := x"4209";
    tmp(13306) := x"4a6b";
    tmp(13307) := x"5acd";
    tmp(13308) := x"630e";
    tmp(13309) := x"6b2e";
    tmp(13310) := x"734f";
    tmp(13311) := x"8bd1";
    tmp(13312) := x"8c13";
    tmp(13313) := x"9413";
    tmp(13314) := x"9c14";
    tmp(13315) := x"7b2f";
    tmp(13316) := x"830e";
    tmp(13317) := x"b453";
    tmp(13318) := x"b474";
    tmp(13319) := x"9391";
    tmp(13320) := x"ac54";
    tmp(13321) := x"ac14";
    tmp(13322) := x"bc75";
    tmp(13323) := x"dcf7";
    tmp(13324) := x"8a8c";
    tmp(13325) := x"b3f1";
    tmp(13326) := x"932e";
    tmp(13327) := x"4146";
    tmp(13328) := x"20a3";
    tmp(13329) := x"0821";
    tmp(13330) := x"0820";
    tmp(13331) := x"1061";
    tmp(13332) := x"28c3";
    tmp(13333) := x"1882";
    tmp(13334) := x"20a3";
    tmp(13335) := x"4187";
    tmp(13336) := x"6a4a";
    tmp(13337) := x"7aab";
    tmp(13338) := x"51a7";
    tmp(13339) := x"726b";
    tmp(13340) := x"932e";
    tmp(13341) := x"ab90";
    tmp(13342) := x"a3af";
    tmp(13343) := x"c4b3";
    tmp(13344) := x"a3ae";
    tmp(13345) := x"b3ef";
    tmp(13346) := x"dcf3";
    tmp(13347) := x"ff1b";
    tmp(13348) := x"ff39";
    tmp(13349) := x"8ae9";
    tmp(13350) := x"0820";
    tmp(13351) := x"0860";
    tmp(13352) := x"08a0";
    tmp(13353) := x"10c0";
    tmp(13354) := x"1100";
    tmp(13355) := x"1940";
    tmp(13356) := x"3200";
    tmp(13357) := x"2a40";
    tmp(13358) := x"08c0";
    tmp(13359) := x"0080";
    tmp(13360) := x"0880";
    tmp(13361) := x"0880";
    tmp(13362) := x"0860";
    tmp(13363) := x"0860";
    tmp(13364) := x"0860";
    tmp(13365) := x"0860";
    tmp(13366) := x"0040";
    tmp(13367) := x"0040";
    tmp(13368) := x"0840";
    tmp(13369) := x"0840";
    tmp(13370) := x"0840";
    tmp(13371) := x"0840";
    tmp(13372) := x"0840";
    tmp(13373) := x"0840";
    tmp(13374) := x"0840";
    tmp(13375) := x"0840";
    tmp(13376) := x"0840";
    tmp(13377) := x"0840";
    tmp(13378) := x"0840";
    tmp(13379) := x"0840";
    tmp(13380) := x"0840";
    tmp(13381) := x"0840";
    tmp(13382) := x"0840";
    tmp(13383) := x"0840";
    tmp(13384) := x"0840";
    tmp(13385) := x"0840";
    tmp(13386) := x"0860";
    tmp(13387) := x"0860";
    tmp(13388) := x"0860";
    tmp(13389) := x"0860";
    tmp(13390) := x"0860";
    tmp(13391) := x"0860";
    tmp(13392) := x"0860";
    tmp(13393) := x"0060";
    tmp(13394) := x"0860";
    tmp(13395) := x"0060";
    tmp(13396) := x"0060";
    tmp(13397) := x"0000";
    tmp(13398) := x"0000";
    tmp(13399) := x"0000";
    tmp(13400) := x"0000";
    tmp(13401) := x"0000";
    tmp(13402) := x"0000";
    tmp(13403) := x"0000";
    tmp(13404) := x"0000";
    tmp(13405) := x"0000";
    tmp(13406) := x"0000";
    tmp(13407) := x"0000";
    tmp(13408) := x"0000";
    tmp(13409) := x"0000";
    tmp(13410) := x"0000";
    tmp(13411) := x"0000";
    tmp(13412) := x"0000";
    tmp(13413) := x"0000";
    tmp(13414) := x"0000";
    tmp(13415) := x"0000";
    tmp(13416) := x"0000";
    tmp(13417) := x"0000";
    tmp(13418) := x"0000";
    tmp(13419) := x"0000";
    tmp(13420) := x"0000";
    tmp(13421) := x"0000";
    tmp(13422) := x"0000";
    tmp(13423) := x"0000";
    tmp(13424) := x"0000";
    tmp(13425) := x"0000";
    tmp(13426) := x"0000";
    tmp(13427) := x"0000";
    tmp(13428) := x"0000";
    tmp(13429) := x"0000";
    tmp(13430) := x"0000";
    tmp(13431) := x"0000";
    tmp(13432) := x"0000";
    tmp(13433) := x"0000";
    tmp(13434) := x"0000";
    tmp(13435) := x"0000";
    tmp(13436) := x"0000";
    tmp(13437) := x"0000";
    tmp(13438) := x"0020";
    tmp(13439) := x"0000";
    tmp(13440) := x"1040";
    tmp(13441) := x"9aa0";
    tmp(13442) := x"9280";
    tmp(13443) := x"9260";
    tmp(13444) := x"8a60";
    tmp(13445) := x"8240";
    tmp(13446) := x"8220";
    tmp(13447) := x"8a40";
    tmp(13448) := x"9240";
    tmp(13449) := x"9a80";
    tmp(13450) := x"a2c0";
    tmp(13451) := x"a2c0";
    tmp(13452) := x"aac0";
    tmp(13453) := x"9a80";
    tmp(13454) := x"aac0";
    tmp(13455) := x"a280";
    tmp(13456) := x"b2a0";
    tmp(13457) := x"b2c0";
    tmp(13458) := x"aa80";
    tmp(13459) := x"b2a0";
    tmp(13460) := x"aa80";
    tmp(13461) := x"aa80";
    tmp(13462) := x"b2a0";
    tmp(13463) := x"bac0";
    tmp(13464) := x"aa80";
    tmp(13465) := x"a260";
    tmp(13466) := x"a260";
    tmp(13467) := x"a260";
    tmp(13468) := x"9a60";
    tmp(13469) := x"9a80";
    tmp(13470) := x"a260";
    tmp(13471) := x"9a60";
    tmp(13472) := x"a260";
    tmp(13473) := x"a280";
    tmp(13474) := x"aaa0";
    tmp(13475) := x"aaa0";
    tmp(13476) := x"aaa0";
    tmp(13477) := x"aac0";
    tmp(13478) := x"b2e0";
    tmp(13479) := x"bb00";
    tmp(13480) := x"b2c0";
    tmp(13481) := x"b2c0";
    tmp(13482) := x"a2a0";
    tmp(13483) := x"aa80";
    tmp(13484) := x"b2c0";
    tmp(13485) := x"d360";
    tmp(13486) := x"c300";
    tmp(13487) := x"b2a0";
    tmp(13488) := x"bac0";
    tmp(13489) := x"b2a0";
    tmp(13490) := x"b2c0";
    tmp(13491) := x"bae0";
    tmp(13492) := x"bac0";
    tmp(13493) := x"bae0";
    tmp(13494) := x"bac0";
    tmp(13495) := x"b2c0";
    tmp(13496) := x"b2c0";
    tmp(13497) := x"bb00";
    tmp(13498) := x"bb00";
    tmp(13499) := x"bb00";
    tmp(13500) := x"bb20";
    tmp(13501) := x"bb20";
    tmp(13502) := x"bb20";
    tmp(13503) := x"b320";
    tmp(13504) := x"b320";
    tmp(13505) := x"aac0";
    tmp(13506) := x"aac0";
    tmp(13507) := x"a2a0";
    tmp(13508) := x"aaa0";
    tmp(13509) := x"aac0";
    tmp(13510) := x"a280";
    tmp(13511) := x"8200";
    tmp(13512) := x"5980";
    tmp(13513) := x"30e0";
    tmp(13514) := x"1060";
    tmp(13515) := x"0820";
    tmp(13516) := x"0000";
    tmp(13517) := x"0000";
    tmp(13518) := x"0000";
    tmp(13519) := x"0000";
    tmp(13520) := x"0000";
    tmp(13521) := x"0000";
    tmp(13522) := x"0000";
    tmp(13523) := x"0000";
    tmp(13524) := x"0000";
    tmp(13525) := x"0000";
    tmp(13526) := x"0000";
    tmp(13527) := x"0000";
    tmp(13528) := x"0000";
    tmp(13529) := x"0000";
    tmp(13530) := x"0000";
    tmp(13531) := x"0000";
    tmp(13532) := x"0000";
    tmp(13533) := x"0000";
    tmp(13534) := x"0000";
    tmp(13535) := x"0000";
    tmp(13536) := x"0000";
    tmp(13537) := x"0000";
    tmp(13538) := x"1061";
    tmp(13539) := x"3966";
    tmp(13540) := x"4187";
    tmp(13541) := x"49c9";
    tmp(13542) := x"5a4a";
    tmp(13543) := x"6aad";
    tmp(13544) := x"6acd";
    tmp(13545) := x"7b70";
    tmp(13546) := x"83b2";
    tmp(13547) := x"8bd3";
    tmp(13548) := x"8b92";
    tmp(13549) := x"834f";
    tmp(13550) := x"9390";
    tmp(13551) := x"9bb1";
    tmp(13552) := x"b496";
    tmp(13553) := x"ac55";
    tmp(13554) := x"8b2f";
    tmp(13555) := x"a3d2";
    tmp(13556) := x"cd17";
    tmp(13557) := x"a3f3";
    tmp(13558) := x"9371";
    tmp(13559) := x"ac13";
    tmp(13560) := x"b455";
    tmp(13561) := x"82cd";
    tmp(13562) := x"ccf5";
    tmp(13563) := x"dd78";
    tmp(13564) := x"724a";
    tmp(13565) := x"4166";
    tmp(13566) := x"0820";
    tmp(13567) := x"0000";
    tmp(13568) := x"0000";
    tmp(13569) := x"1061";
    tmp(13570) := x"72ea";
    tmp(13571) := x"49e7";
    tmp(13572) := x"1861";
    tmp(13573) := x"4185";
    tmp(13574) := x"4165";
    tmp(13575) := x"5a08";
    tmp(13576) := x"51a7";
    tmp(13577) := x"51a7";
    tmp(13578) := x"a3cf";
    tmp(13579) := x"59c8";
    tmp(13580) := x"6a09";
    tmp(13581) := x"ab8f";
    tmp(13582) := x"a36f";
    tmp(13583) := x"a3b0";
    tmp(13584) := x"abaf";
    tmp(13585) := x"e5b5";
    tmp(13586) := x"edd5";
    tmp(13587) := x"edd5";
    tmp(13588) := x"4985";
    tmp(13589) := x"0840";
    tmp(13590) := x"0840";
    tmp(13591) := x"0880";
    tmp(13592) := x"08c0";
    tmp(13593) := x"10e0";
    tmp(13594) := x"1920";
    tmp(13595) := x"2160";
    tmp(13596) := x"3200";
    tmp(13597) := x"3240";
    tmp(13598) := x"08e0";
    tmp(13599) := x"0080";
    tmp(13600) := x"08a0";
    tmp(13601) := x"0880";
    tmp(13602) := x"0880";
    tmp(13603) := x"0880";
    tmp(13604) := x"0880";
    tmp(13605) := x"0060";
    tmp(13606) := x"0860";
    tmp(13607) := x"0860";
    tmp(13608) := x"0840";
    tmp(13609) := x"0840";
    tmp(13610) := x"0840";
    tmp(13611) := x"0840";
    tmp(13612) := x"0840";
    tmp(13613) := x"0840";
    tmp(13614) := x"0840";
    tmp(13615) := x"0840";
    tmp(13616) := x"0840";
    tmp(13617) := x"0840";
    tmp(13618) := x"0840";
    tmp(13619) := x"0840";
    tmp(13620) := x"0840";
    tmp(13621) := x"0840";
    tmp(13622) := x"0840";
    tmp(13623) := x"0840";
    tmp(13624) := x"0840";
    tmp(13625) := x"0840";
    tmp(13626) := x"0840";
    tmp(13627) := x"0840";
    tmp(13628) := x"0840";
    tmp(13629) := x"0840";
    tmp(13630) := x"0840";
    tmp(13631) := x"0860";
    tmp(13632) := x"0860";
    tmp(13633) := x"0860";
    tmp(13634) := x"0060";
    tmp(13635) := x"0060";
    tmp(13636) := x"0060";
    tmp(13637) := x"0000";
    tmp(13638) := x"0000";
    tmp(13639) := x"0000";
    tmp(13640) := x"0000";
    tmp(13641) := x"0000";
    tmp(13642) := x"0000";
    tmp(13643) := x"0000";
    tmp(13644) := x"0000";
    tmp(13645) := x"0000";
    tmp(13646) := x"0000";
    tmp(13647) := x"0000";
    tmp(13648) := x"0000";
    tmp(13649) := x"0000";
    tmp(13650) := x"0000";
    tmp(13651) := x"0000";
    tmp(13652) := x"0000";
    tmp(13653) := x"0000";
    tmp(13654) := x"0000";
    tmp(13655) := x"0000";
    tmp(13656) := x"0000";
    tmp(13657) := x"0000";
    tmp(13658) := x"0000";
    tmp(13659) := x"0000";
    tmp(13660) := x"0000";
    tmp(13661) := x"0000";
    tmp(13662) := x"0000";
    tmp(13663) := x"0000";
    tmp(13664) := x"0000";
    tmp(13665) := x"0000";
    tmp(13666) := x"0000";
    tmp(13667) := x"0000";
    tmp(13668) := x"0000";
    tmp(13669) := x"0000";
    tmp(13670) := x"0000";
    tmp(13671) := x"0000";
    tmp(13672) := x"0000";
    tmp(13673) := x"0000";
    tmp(13674) := x"0000";
    tmp(13675) := x"0000";
    tmp(13676) := x"0000";
    tmp(13677) := x"0020";
    tmp(13678) := x"0000";
    tmp(13679) := x"0020";
    tmp(13680) := x"1040";
    tmp(13681) := x"b2e0";
    tmp(13682) := x"aac0";
    tmp(13683) := x"aac0";
    tmp(13684) := x"aac0";
    tmp(13685) := x"a280";
    tmp(13686) := x"a2a0";
    tmp(13687) := x"aac0";
    tmp(13688) := x"b2a0";
    tmp(13689) := x"aaa0";
    tmp(13690) := x"aac0";
    tmp(13691) := x"aac0";
    tmp(13692) := x"aac0";
    tmp(13693) := x"aac0";
    tmp(13694) := x"b2e0";
    tmp(13695) := x"bae0";
    tmp(13696) := x"bac0";
    tmp(13697) := x"b2a0";
    tmp(13698) := x"b2c0";
    tmp(13699) := x"b2a0";
    tmp(13700) := x"aa80";
    tmp(13701) := x"b2a0";
    tmp(13702) := x"b2a0";
    tmp(13703) := x"aa80";
    tmp(13704) := x"aa80";
    tmp(13705) := x"aa80";
    tmp(13706) := x"a260";
    tmp(13707) := x"9a40";
    tmp(13708) := x"9240";
    tmp(13709) := x"9240";
    tmp(13710) := x"9240";
    tmp(13711) := x"9a60";
    tmp(13712) := x"9a60";
    tmp(13713) := x"aac0";
    tmp(13714) := x"aac0";
    tmp(13715) := x"aaa0";
    tmp(13716) := x"aaa0";
    tmp(13717) := x"aac0";
    tmp(13718) := x"b2c0";
    tmp(13719) := x"aaa0";
    tmp(13720) := x"aa80";
    tmp(13721) := x"a280";
    tmp(13722) := x"a280";
    tmp(13723) := x"aa80";
    tmp(13724) := x"b2c0";
    tmp(13725) := x"b2e0";
    tmp(13726) := x"bb00";
    tmp(13727) := x"b2c0";
    tmp(13728) := x"aa80";
    tmp(13729) := x"b2c0";
    tmp(13730) := x"bae0";
    tmp(13731) := x"b2c0";
    tmp(13732) := x"aa80";
    tmp(13733) := x"aa80";
    tmp(13734) := x"a280";
    tmp(13735) := x"a260";
    tmp(13736) := x"a260";
    tmp(13737) := x"b2c0";
    tmp(13738) := x"b2c0";
    tmp(13739) := x"b2a0";
    tmp(13740) := x"b2a0";
    tmp(13741) := x"b2e0";
    tmp(13742) := x"b300";
    tmp(13743) := x"bb20";
    tmp(13744) := x"b2e0";
    tmp(13745) := x"aaa0";
    tmp(13746) := x"a280";
    tmp(13747) := x"aaa0";
    tmp(13748) := x"aaa0";
    tmp(13749) := x"aac0";
    tmp(13750) := x"a280";
    tmp(13751) := x"8220";
    tmp(13752) := x"5180";
    tmp(13753) := x"28c0";
    tmp(13754) := x"0840";
    tmp(13755) := x"0020";
    tmp(13756) := x"0000";
    tmp(13757) := x"0000";
    tmp(13758) := x"0000";
    tmp(13759) := x"0020";
    tmp(13760) := x"0020";
    tmp(13761) := x"0000";
    tmp(13762) := x"0000";
    tmp(13763) := x"0000";
    tmp(13764) := x"0000";
    tmp(13765) := x"0000";
    tmp(13766) := x"0000";
    tmp(13767) := x"0000";
    tmp(13768) := x"0000";
    tmp(13769) := x"0000";
    tmp(13770) := x"0000";
    tmp(13771) := x"0000";
    tmp(13772) := x"0000";
    tmp(13773) := x"0000";
    tmp(13774) := x"0000";
    tmp(13775) := x"0000";
    tmp(13776) := x"0000";
    tmp(13777) := x"0000";
    tmp(13778) := x"20a2";
    tmp(13779) := x"4987";
    tmp(13780) := x"4188";
    tmp(13781) := x"49a9";
    tmp(13782) := x"5a4b";
    tmp(13783) := x"5a4c";
    tmp(13784) := x"49c9";
    tmp(13785) := x"6a8d";
    tmp(13786) := x"8b92";
    tmp(13787) := x"8372";
    tmp(13788) := x"8372";
    tmp(13789) := x"8b71";
    tmp(13790) := x"8b71";
    tmp(13791) := x"ac54";
    tmp(13792) := x"cd79";
    tmp(13793) := x"bcf7";
    tmp(13794) := x"b453";
    tmp(13795) := x"cd38";
    tmp(13796) := x"ac56";
    tmp(13797) := x"93b3";
    tmp(13798) := x"bc97";
    tmp(13799) := x"b456";
    tmp(13800) := x"9371";
    tmp(13801) := x"9b6e";
    tmp(13802) := x"fedc";
    tmp(13803) := x"930d";
    tmp(13804) := x"3925";
    tmp(13805) := x"20c3";
    tmp(13806) := x"0820";
    tmp(13807) := x"0820";
    tmp(13808) := x"3944";
    tmp(13809) := x"72a9";
    tmp(13810) := x"6a6a";
    tmp(13811) := x"0820";
    tmp(13812) := x"3124";
    tmp(13813) := x"51e7";
    tmp(13814) := x"3924";
    tmp(13815) := x"51e8";
    tmp(13816) := x"4145";
    tmp(13817) := x"4165";
    tmp(13818) := x"edf9";
    tmp(13819) := x"ccf5";
    tmp(13820) := x"92ec";
    tmp(13821) := x"7229";
    tmp(13822) := x"6a08";
    tmp(13823) := x"9b0d";
    tmp(13824) := x"92cb";
    tmp(13825) := x"ccf2";
    tmp(13826) := x"6a68";
    tmp(13827) := x"1881";
    tmp(13828) := x"0820";
    tmp(13829) := x"0860";
    tmp(13830) := x"0880";
    tmp(13831) := x"10c0";
    tmp(13832) := x"10e0";
    tmp(13833) := x"10e0";
    tmp(13834) := x"1900";
    tmp(13835) := x"2160";
    tmp(13836) := x"29e0";
    tmp(13837) := x"3ac1";
    tmp(13838) := x"1140";
    tmp(13839) := x"00a0";
    tmp(13840) := x"08a0";
    tmp(13841) := x"08a0";
    tmp(13842) := x"0880";
    tmp(13843) := x"0880";
    tmp(13844) := x"0880";
    tmp(13845) := x"0880";
    tmp(13846) := x"0860";
    tmp(13847) := x"0860";
    tmp(13848) := x"0860";
    tmp(13849) := x"0860";
    tmp(13850) := x"0840";
    tmp(13851) := x"0840";
    tmp(13852) := x"0840";
    tmp(13853) := x"0840";
    tmp(13854) := x"0840";
    tmp(13855) := x"0840";
    tmp(13856) := x"0840";
    tmp(13857) := x"0840";
    tmp(13858) := x"0840";
    tmp(13859) := x"0840";
    tmp(13860) := x"0820";
    tmp(13861) := x"0820";
    tmp(13862) := x"0840";
    tmp(13863) := x"0840";
    tmp(13864) := x"0840";
    tmp(13865) := x"0840";
    tmp(13866) := x"0840";
    tmp(13867) := x"0840";
    tmp(13868) := x"0840";
    tmp(13869) := x"0840";
    tmp(13870) := x"0840";
    tmp(13871) := x"0840";
    tmp(13872) := x"0840";
    tmp(13873) := x"0840";
    tmp(13874) := x"0040";
    tmp(13875) := x"0040";
    tmp(13876) := x"0060";
    tmp(13877) := x"0000";
    tmp(13878) := x"0000";
    tmp(13879) := x"0000";
    tmp(13880) := x"0000";
    tmp(13881) := x"0000";
    tmp(13882) := x"0000";
    tmp(13883) := x"0000";
    tmp(13884) := x"0000";
    tmp(13885) := x"0000";
    tmp(13886) := x"0000";
    tmp(13887) := x"0000";
    tmp(13888) := x"0000";
    tmp(13889) := x"0000";
    tmp(13890) := x"0000";
    tmp(13891) := x"0000";
    tmp(13892) := x"0000";
    tmp(13893) := x"0000";
    tmp(13894) := x"0000";
    tmp(13895) := x"0000";
    tmp(13896) := x"0000";
    tmp(13897) := x"0000";
    tmp(13898) := x"0000";
    tmp(13899) := x"0000";
    tmp(13900) := x"0000";
    tmp(13901) := x"0000";
    tmp(13902) := x"0000";
    tmp(13903) := x"0000";
    tmp(13904) := x"0000";
    tmp(13905) := x"0000";
    tmp(13906) := x"0000";
    tmp(13907) := x"0000";
    tmp(13908) := x"0000";
    tmp(13909) := x"0000";
    tmp(13910) := x"0000";
    tmp(13911) := x"0000";
    tmp(13912) := x"0000";
    tmp(13913) := x"0000";
    tmp(13914) := x"0000";
    tmp(13915) := x"0000";
    tmp(13916) := x"0000";
    tmp(13917) := x"0000";
    tmp(13918) := x"0020";
    tmp(13919) := x"0000";
    tmp(13920) := x"1040";
    tmp(13921) := x"c340";
    tmp(13922) := x"b300";
    tmp(13923) := x"bb40";
    tmp(13924) := x"bb40";
    tmp(13925) := x"c320";
    tmp(13926) := x"bb20";
    tmp(13927) := x"bb20";
    tmp(13928) := x"c320";
    tmp(13929) := x"c320";
    tmp(13930) := x"c300";
    tmp(13931) := x"bb00";
    tmp(13932) := x"bb00";
    tmp(13933) := x"b2c0";
    tmp(13934) := x"b2c0";
    tmp(13935) := x"c300";
    tmp(13936) := x"c300";
    tmp(13937) := x"bac0";
    tmp(13938) := x"bac0";
    tmp(13939) := x"c2e0";
    tmp(13940) := x"baa0";
    tmp(13941) := x"baa0";
    tmp(13942) := x"b2a0";
    tmp(13943) := x"aa80";
    tmp(13944) := x"a240";
    tmp(13945) := x"a240";
    tmp(13946) := x"9a40";
    tmp(13947) := x"9240";
    tmp(13948) := x"9240";
    tmp(13949) := x"9220";
    tmp(13950) := x"9240";
    tmp(13951) := x"9a40";
    tmp(13952) := x"9a60";
    tmp(13953) := x"a280";
    tmp(13954) := x"aac0";
    tmp(13955) := x"b2c0";
    tmp(13956) := x"aac0";
    tmp(13957) := x"aac0";
    tmp(13958) := x"aaa0";
    tmp(13959) := x"a280";
    tmp(13960) := x"9a60";
    tmp(13961) := x"9a60";
    tmp(13962) := x"a280";
    tmp(13963) := x"aaa0";
    tmp(13964) := x"aac0";
    tmp(13965) := x"aaa0";
    tmp(13966) := x"aa80";
    tmp(13967) := x"aaa0";
    tmp(13968) := x"aaa0";
    tmp(13969) := x"b2c0";
    tmp(13970) := x"b2c0";
    tmp(13971) := x"aaa0";
    tmp(13972) := x"aa80";
    tmp(13973) := x"a280";
    tmp(13974) := x"a260";
    tmp(13975) := x"a240";
    tmp(13976) := x"9200";
    tmp(13977) := x"81c0";
    tmp(13978) := x"89c0";
    tmp(13979) := x"a240";
    tmp(13980) := x"a260";
    tmp(13981) := x"b2c0";
    tmp(13982) := x"b2c0";
    tmp(13983) := x"b2c0";
    tmp(13984) := x"b2c0";
    tmp(13985) := x"b2c0";
    tmp(13986) := x"b2e0";
    tmp(13987) := x"b2e0";
    tmp(13988) := x"b2c0";
    tmp(13989) := x"aaa0";
    tmp(13990) := x"9a60";
    tmp(13991) := x"7a00";
    tmp(13992) := x"4140";
    tmp(13993) := x"1880";
    tmp(13994) := x"0840";
    tmp(13995) := x"0020";
    tmp(13996) := x"0000";
    tmp(13997) := x"0000";
    tmp(13998) := x"0000";
    tmp(13999) := x"0020";
    tmp(14000) := x"0020";
    tmp(14001) := x"0000";
    tmp(14002) := x"0000";
    tmp(14003) := x"0000";
    tmp(14004) := x"0000";
    tmp(14005) := x"0000";
    tmp(14006) := x"0000";
    tmp(14007) := x"0000";
    tmp(14008) := x"0000";
    tmp(14009) := x"0000";
    tmp(14010) := x"0000";
    tmp(14011) := x"0000";
    tmp(14012) := x"0000";
    tmp(14013) := x"0000";
    tmp(14014) := x"0000";
    tmp(14015) := x"0000";
    tmp(14016) := x"0000";
    tmp(14017) := x"0820";
    tmp(14018) := x"3925";
    tmp(14019) := x"4187";
    tmp(14020) := x"5a2b";
    tmp(14021) := x"6a8d";
    tmp(14022) := x"522b";
    tmp(14023) := x"522b";
    tmp(14024) := x"6aad";
    tmp(14025) := x"72ef";
    tmp(14026) := x"7b51";
    tmp(14027) := x"93b3";
    tmp(14028) := x"8bb2";
    tmp(14029) := x"9c54";
    tmp(14030) := x"bcf8";
    tmp(14031) := x"c558";
    tmp(14032) := x"d5b9";
    tmp(14033) := x"e65c";
    tmp(14034) := x"f69e";
    tmp(14035) := x"c55a";
    tmp(14036) := x"bcf8";
    tmp(14037) := x"e5fd";
    tmp(14038) := x"9bf4";
    tmp(14039) := x"ccf9";
    tmp(14040) := x"9b70";
    tmp(14041) := x"d535";
    tmp(14042) := x"edf9";
    tmp(14043) := x"59e8";
    tmp(14044) := x"0820";
    tmp(14045) := x"0000";
    tmp(14046) := x"0000";
    tmp(14047) := x"1041";
    tmp(14048) := x"5a08";
    tmp(14049) := x"6229";
    tmp(14050) := x"1041";
    tmp(14051) := x"1061";
    tmp(14052) := x"ac50";
    tmp(14053) := x"1882";
    tmp(14054) := x"4165";
    tmp(14055) := x"20a2";
    tmp(14056) := x"6248";
    tmp(14057) := x"3104";
    tmp(14058) := x"ccd5";
    tmp(14059) := x"d517";
    tmp(14060) := x"fdf9";
    tmp(14061) := x"9b4d";
    tmp(14062) := x"7249";
    tmp(14063) := x"828a";
    tmp(14064) := x"ab8d";
    tmp(14065) := x"59e7";
    tmp(14066) := x"0820";
    tmp(14067) := x"0840";
    tmp(14068) := x"0880";
    tmp(14069) := x"0880";
    tmp(14070) := x"0880";
    tmp(14071) := x"10c0";
    tmp(14072) := x"10e0";
    tmp(14073) := x"10e0";
    tmp(14074) := x"1920";
    tmp(14075) := x"2180";
    tmp(14076) := x"29e0";
    tmp(14077) := x"3ac1";
    tmp(14078) := x"1160";
    tmp(14079) := x"08a0";
    tmp(14080) := x"08c0";
    tmp(14081) := x"08a0";
    tmp(14082) := x"08a0";
    tmp(14083) := x"08a0";
    tmp(14084) := x"08a0";
    tmp(14085) := x"0880";
    tmp(14086) := x"0880";
    tmp(14087) := x"0880";
    tmp(14088) := x"0860";
    tmp(14089) := x"0860";
    tmp(14090) := x"0860";
    tmp(14091) := x"0860";
    tmp(14092) := x"0860";
    tmp(14093) := x"0840";
    tmp(14094) := x"0840";
    tmp(14095) := x"0840";
    tmp(14096) := x"0840";
    tmp(14097) := x"0840";
    tmp(14098) := x"0840";
    tmp(14099) := x"0840";
    tmp(14100) := x"0820";
    tmp(14101) := x"0820";
    tmp(14102) := x"0820";
    tmp(14103) := x"0820";
    tmp(14104) := x"0820";
    tmp(14105) := x"0820";
    tmp(14106) := x"0820";
    tmp(14107) := x"0820";
    tmp(14108) := x"0840";
    tmp(14109) := x"0840";
    tmp(14110) := x"0840";
    tmp(14111) := x"0840";
    tmp(14112) := x"0840";
    tmp(14113) := x"0840";
    tmp(14114) := x"0840";
    tmp(14115) := x"0040";
    tmp(14116) := x"0040";
    tmp(14117) := x"0000";
    tmp(14118) := x"0000";
    tmp(14119) := x"0000";
    tmp(14120) := x"0000";
    tmp(14121) := x"0000";
    tmp(14122) := x"0000";
    tmp(14123) := x"0000";
    tmp(14124) := x"0000";
    tmp(14125) := x"0000";
    tmp(14126) := x"0000";
    tmp(14127) := x"0000";
    tmp(14128) := x"0000";
    tmp(14129) := x"0000";
    tmp(14130) := x"0000";
    tmp(14131) := x"0000";
    tmp(14132) := x"0000";
    tmp(14133) := x"0000";
    tmp(14134) := x"0000";
    tmp(14135) := x"0000";
    tmp(14136) := x"0000";
    tmp(14137) := x"0000";
    tmp(14138) := x"0000";
    tmp(14139) := x"0000";
    tmp(14140) := x"0000";
    tmp(14141) := x"0000";
    tmp(14142) := x"0000";
    tmp(14143) := x"0000";
    tmp(14144) := x"0000";
    tmp(14145) := x"0000";
    tmp(14146) := x"0000";
    tmp(14147) := x"0000";
    tmp(14148) := x"0000";
    tmp(14149) := x"0000";
    tmp(14150) := x"0000";
    tmp(14151) := x"0000";
    tmp(14152) := x"0000";
    tmp(14153) := x"0000";
    tmp(14154) := x"0000";
    tmp(14155) := x"0000";
    tmp(14156) := x"0000";
    tmp(14157) := x"0020";
    tmp(14158) := x"0020";
    tmp(14159) := x"0020";
    tmp(14160) := x"1040";
    tmp(14161) := x"bb20";
    tmp(14162) := x"b2e0";
    tmp(14163) := x"c340";
    tmp(14164) := x"cb40";
    tmp(14165) := x"d380";
    tmp(14166) := x"d3a0";
    tmp(14167) := x"dba0";
    tmp(14168) := x"d380";
    tmp(14169) := x"cb60";
    tmp(14170) := x"cb60";
    tmp(14171) := x"c340";
    tmp(14172) := x"cb40";
    tmp(14173) := x"bb20";
    tmp(14174) := x"c340";
    tmp(14175) := x"bb20";
    tmp(14176) := x"cb20";
    tmp(14177) := x"c2c0";
    tmp(14178) := x"bac0";
    tmp(14179) := x"c2e0";
    tmp(14180) := x"c2c0";
    tmp(14181) := x"c2c0";
    tmp(14182) := x"bac0";
    tmp(14183) := x"aa60";
    tmp(14184) := x"9a20";
    tmp(14185) := x"9220";
    tmp(14186) := x"9220";
    tmp(14187) := x"8a00";
    tmp(14188) := x"9200";
    tmp(14189) := x"8a00";
    tmp(14190) := x"9220";
    tmp(14191) := x"9200";
    tmp(14192) := x"9a40";
    tmp(14193) := x"a260";
    tmp(14194) := x"aac0";
    tmp(14195) := x"b2e0";
    tmp(14196) := x"aac0";
    tmp(14197) := x"b2c0";
    tmp(14198) := x"aaa0";
    tmp(14199) := x"a280";
    tmp(14200) := x"9a60";
    tmp(14201) := x"9a60";
    tmp(14202) := x"a280";
    tmp(14203) := x"aaa0";
    tmp(14204) := x"aaa0";
    tmp(14205) := x"a2a0";
    tmp(14206) := x"a280";
    tmp(14207) := x"b2a0";
    tmp(14208) := x"aa80";
    tmp(14209) := x"aaa0";
    tmp(14210) := x"aaa0";
    tmp(14211) := x"a280";
    tmp(14212) := x"a260";
    tmp(14213) := x"a280";
    tmp(14214) := x"a260";
    tmp(14215) := x"a240";
    tmp(14216) := x"9a20";
    tmp(14217) := x"89e0";
    tmp(14218) := x"79a0";
    tmp(14219) := x"7180";
    tmp(14220) := x"79a0";
    tmp(14221) := x"89c0";
    tmp(14222) := x"89e0";
    tmp(14223) := x"9220";
    tmp(14224) := x"9240";
    tmp(14225) := x"9a60";
    tmp(14226) := x"aac0";
    tmp(14227) := x"aac0";
    tmp(14228) := x"aac0";
    tmp(14229) := x"aac0";
    tmp(14230) := x"9a60";
    tmp(14231) := x"71e0";
    tmp(14232) := x"3920";
    tmp(14233) := x"1880";
    tmp(14234) := x"0820";
    tmp(14235) := x"0020";
    tmp(14236) := x"0000";
    tmp(14237) := x"0000";
    tmp(14238) := x"0000";
    tmp(14239) := x"0020";
    tmp(14240) := x"0000";
    tmp(14241) := x"0000";
    tmp(14242) := x"0000";
    tmp(14243) := x"0000";
    tmp(14244) := x"0000";
    tmp(14245) := x"0000";
    tmp(14246) := x"0000";
    tmp(14247) := x"0000";
    tmp(14248) := x"0000";
    tmp(14249) := x"0000";
    tmp(14250) := x"0000";
    tmp(14251) := x"0000";
    tmp(14252) := x"0000";
    tmp(14253) := x"0000";
    tmp(14254) := x"0000";
    tmp(14255) := x"0000";
    tmp(14256) := x"0000";
    tmp(14257) := x"1041";
    tmp(14258) := x"49a6";
    tmp(14259) := x"6a8b";
    tmp(14260) := x"72ee";
    tmp(14261) := x"6acf";
    tmp(14262) := x"6a8d";
    tmp(14263) := x"6aad";
    tmp(14264) := x"6a8d";
    tmp(14265) := x"8351";
    tmp(14266) := x"93d3";
    tmp(14267) := x"93d2";
    tmp(14268) := x"ac76";
    tmp(14269) := x"c518";
    tmp(14270) := x"cd39";
    tmp(14271) := x"cd7a";
    tmp(14272) := x"e69c";
    tmp(14273) := x"f6ff";
    tmp(14274) := x"ee3d";
    tmp(14275) := x"dd7a";
    tmp(14276) := x"ee5e";
    tmp(14277) := x"b4d8";
    tmp(14278) := x"ddbb";
    tmp(14279) := x"b414";
    tmp(14280) := x"c4f5";
    tmp(14281) := x"ff5d";
    tmp(14282) := x"e5f9";
    tmp(14283) := x"3125";
    tmp(14284) := x"0841";
    tmp(14285) := x"0820";
    tmp(14286) := x"1041";
    tmp(14287) := x"728a";
    tmp(14288) := x"832c";
    tmp(14289) := x"0841";
    tmp(14290) := x"1881";
    tmp(14291) := x"832b";
    tmp(14292) := x"6249";
    tmp(14293) := x"0821";
    tmp(14294) := x"728a";
    tmp(14295) := x"5a08";
    tmp(14296) := x"6a6a";
    tmp(14297) := x"20a3";
    tmp(14298) := x"728b";
    tmp(14299) := x"932e";
    tmp(14300) := x"f5d9";
    tmp(14301) := x"ed76";
    tmp(14302) := x"d534";
    tmp(14303) := x"b490";
    tmp(14304) := x"dd33";
    tmp(14305) := x"20c2";
    tmp(14306) := x"0840";
    tmp(14307) := x"08a0";
    tmp(14308) := x"08c0";
    tmp(14309) := x"08a0";
    tmp(14310) := x"10a0";
    tmp(14311) := x"10e0";
    tmp(14312) := x"1120";
    tmp(14313) := x"10e0";
    tmp(14314) := x"1940";
    tmp(14315) := x"2180";
    tmp(14316) := x"2180";
    tmp(14317) := x"3260";
    tmp(14318) := x"1160";
    tmp(14319) := x"08a0";
    tmp(14320) := x"08c0";
    tmp(14321) := x"08a0";
    tmp(14322) := x"08a0";
    tmp(14323) := x"08a0";
    tmp(14324) := x"08a0";
    tmp(14325) := x"08a0";
    tmp(14326) := x"08a0";
    tmp(14327) := x"0880";
    tmp(14328) := x"0880";
    tmp(14329) := x"0880";
    tmp(14330) := x"0880";
    tmp(14331) := x"0860";
    tmp(14332) := x"0860";
    tmp(14333) := x"0860";
    tmp(14334) := x"0860";
    tmp(14335) := x"0840";
    tmp(14336) := x"0840";
    tmp(14337) := x"0840";
    tmp(14338) := x"0840";
    tmp(14339) := x"0840";
    tmp(14340) := x"0820";
    tmp(14341) := x"0820";
    tmp(14342) := x"0820";
    tmp(14343) := x"0820";
    tmp(14344) := x"0820";
    tmp(14345) := x"0820";
    tmp(14346) := x"0820";
    tmp(14347) := x"0820";
    tmp(14348) := x"0820";
    tmp(14349) := x"0820";
    tmp(14350) := x"0820";
    tmp(14351) := x"0820";
    tmp(14352) := x"0840";
    tmp(14353) := x"0840";
    tmp(14354) := x"0840";
    tmp(14355) := x"0840";
    tmp(14356) := x"0040";
    tmp(14357) := x"0000";
    tmp(14358) := x"0000";
    tmp(14359) := x"0000";
    tmp(14360) := x"0000";
    tmp(14361) := x"0000";
    tmp(14362) := x"0000";
    tmp(14363) := x"0000";
    tmp(14364) := x"0000";
    tmp(14365) := x"0000";
    tmp(14366) := x"0000";
    tmp(14367) := x"0000";
    tmp(14368) := x"0000";
    tmp(14369) := x"0000";
    tmp(14370) := x"0000";
    tmp(14371) := x"0000";
    tmp(14372) := x"0000";
    tmp(14373) := x"0000";
    tmp(14374) := x"0000";
    tmp(14375) := x"0000";
    tmp(14376) := x"0000";
    tmp(14377) := x"0000";
    tmp(14378) := x"0000";
    tmp(14379) := x"0000";
    tmp(14380) := x"0000";
    tmp(14381) := x"0000";
    tmp(14382) := x"0000";
    tmp(14383) := x"0000";
    tmp(14384) := x"0000";
    tmp(14385) := x"0000";
    tmp(14386) := x"0000";
    tmp(14387) := x"0000";
    tmp(14388) := x"0000";
    tmp(14389) := x"0000";
    tmp(14390) := x"0000";
    tmp(14391) := x"0000";
    tmp(14392) := x"0000";
    tmp(14393) := x"0000";
    tmp(14394) := x"0000";
    tmp(14395) := x"0000";
    tmp(14396) := x"0000";
    tmp(14397) := x"0020";
    tmp(14398) := x"0020";
    tmp(14399) := x"0020";
    tmp(14400) := x"1040";
    tmp(14401) := x"c320";
    tmp(14402) := x"bb00";
    tmp(14403) := x"cb40";
    tmp(14404) := x"cb40";
    tmp(14405) := x"cb60";
    tmp(14406) := x"d3a0";
    tmp(14407) := x"dba0";
    tmp(14408) := x"dba0";
    tmp(14409) := x"d3a0";
    tmp(14410) := x"d3c0";
    tmp(14411) := x"cb80";
    tmp(14412) := x"cb60";
    tmp(14413) := x"cb80";
    tmp(14414) := x"c340";
    tmp(14415) := x"c320";
    tmp(14416) := x"c320";
    tmp(14417) := x"c300";
    tmp(14418) := x"bac0";
    tmp(14419) := x"bac0";
    tmp(14420) := x"c2c0";
    tmp(14421) := x"c2c0";
    tmp(14422) := x"baa0";
    tmp(14423) := x"a260";
    tmp(14424) := x"9a40";
    tmp(14425) := x"9a20";
    tmp(14426) := x"9220";
    tmp(14427) := x"8a20";
    tmp(14428) := x"9220";
    tmp(14429) := x"9200";
    tmp(14430) := x"9200";
    tmp(14431) := x"9a40";
    tmp(14432) := x"aa80";
    tmp(14433) := x"aa80";
    tmp(14434) := x"b2e0";
    tmp(14435) := x"b2e0";
    tmp(14436) := x"aac0";
    tmp(14437) := x"aaa0";
    tmp(14438) := x"aa80";
    tmp(14439) := x"9a60";
    tmp(14440) := x"9a80";
    tmp(14441) := x"9a80";
    tmp(14442) := x"a2a0";
    tmp(14443) := x"aac0";
    tmp(14444) := x"a2a0";
    tmp(14445) := x"a280";
    tmp(14446) := x"a280";
    tmp(14447) := x"aa80";
    tmp(14448) := x"aa80";
    tmp(14449) := x"a260";
    tmp(14450) := x"9a40";
    tmp(14451) := x"9a40";
    tmp(14452) := x"a260";
    tmp(14453) := x"aa60";
    tmp(14454) := x"a260";
    tmp(14455) := x"a220";
    tmp(14456) := x"9a20";
    tmp(14457) := x"9220";
    tmp(14458) := x"9200";
    tmp(14459) := x"81c0";
    tmp(14460) := x"79a0";
    tmp(14461) := x"7180";
    tmp(14462) := x"7160";
    tmp(14463) := x"7160";
    tmp(14464) := x"7180";
    tmp(14465) := x"79c0";
    tmp(14466) := x"8a00";
    tmp(14467) := x"9240";
    tmp(14468) := x"9a80";
    tmp(14469) := x"9a80";
    tmp(14470) := x"8a60";
    tmp(14471) := x"59a0";
    tmp(14472) := x"20c0";
    tmp(14473) := x"1060";
    tmp(14474) := x"0820";
    tmp(14475) := x"0020";
    tmp(14476) := x"0000";
    tmp(14477) := x"0000";
    tmp(14478) := x"0000";
    tmp(14479) := x"0000";
    tmp(14480) := x"0000";
    tmp(14481) := x"0000";
    tmp(14482) := x"0000";
    tmp(14483) := x"0000";
    tmp(14484) := x"0000";
    tmp(14485) := x"0000";
    tmp(14486) := x"0000";
    tmp(14487) := x"0000";
    tmp(14488) := x"0000";
    tmp(14489) := x"0000";
    tmp(14490) := x"0000";
    tmp(14491) := x"0000";
    tmp(14492) := x"0000";
    tmp(14493) := x"0000";
    tmp(14494) := x"0000";
    tmp(14495) := x"0000";
    tmp(14496) := x"0000";
    tmp(14497) := x"1882";
    tmp(14498) := x"6a8a";
    tmp(14499) := x"7b2e";
    tmp(14500) := x"72cd";
    tmp(14501) := x"730f";
    tmp(14502) := x"6a8d";
    tmp(14503) := x"72ad";
    tmp(14504) := x"7ace";
    tmp(14505) := x"8b71";
    tmp(14506) := x"9bd3";
    tmp(14507) := x"b4b6";
    tmp(14508) := x"ac75";
    tmp(14509) := x"ac34";
    tmp(14510) := x"bc95";
    tmp(14511) := x"e63b";
    tmp(14512) := x"ff1f";
    tmp(14513) := x"edbb";
    tmp(14514) := x"e559";
    tmp(14515) := x"fe7d";
    tmp(14516) := x"d59c";
    tmp(14517) := x"bcd7";
    tmp(14518) := x"dd7a";
    tmp(14519) := x"ccd5";
    tmp(14520) := x"ffff";
    tmp(14521) := x"ff1d";
    tmp(14522) := x"8bcf";
    tmp(14523) := x"1041";
    tmp(14524) := x"0000";
    tmp(14525) := x"0020";
    tmp(14526) := x"3104";
    tmp(14527) := x"9bd0";
    tmp(14528) := x"20a2";
    tmp(14529) := x"0820";
    tmp(14530) := x"6269";
    tmp(14531) := x"bc72";
    tmp(14532) := x"1041";
    tmp(14533) := x"20c3";
    tmp(14534) := x"5a29";
    tmp(14535) := x"3945";
    tmp(14536) := x"8b4e";
    tmp(14537) := x"3104";
    tmp(14538) := x"20a3";
    tmp(14539) := x"28c3";
    tmp(14540) := x"8aec";
    tmp(14541) := x"ed97";
    tmp(14542) := x"e535";
    tmp(14543) := x"ee79";
    tmp(14544) := x"cd73";
    tmp(14545) := x"18c1";
    tmp(14546) := x"08a0";
    tmp(14547) := x"08c0";
    tmp(14548) := x"08a0";
    tmp(14549) := x"08a0";
    tmp(14550) := x"10a0";
    tmp(14551) := x"10e0";
    tmp(14552) := x"10e0";
    tmp(14553) := x"1100";
    tmp(14554) := x"2180";
    tmp(14555) := x"2180";
    tmp(14556) := x"21a0";
    tmp(14557) := x"2a20";
    tmp(14558) := x"1140";
    tmp(14559) := x"08a0";
    tmp(14560) := x"08c0";
    tmp(14561) := x"08c0";
    tmp(14562) := x"08c0";
    tmp(14563) := x"08a0";
    tmp(14564) := x"08c0";
    tmp(14565) := x"08c0";
    tmp(14566) := x"08a0";
    tmp(14567) := x"08a0";
    tmp(14568) := x"08a0";
    tmp(14569) := x"08a0";
    tmp(14570) := x"0880";
    tmp(14571) := x"0880";
    tmp(14572) := x"0880";
    tmp(14573) := x"0860";
    tmp(14574) := x"0860";
    tmp(14575) := x"0860";
    tmp(14576) := x"0860";
    tmp(14577) := x"0840";
    tmp(14578) := x"0840";
    tmp(14579) := x"0840";
    tmp(14580) := x"0840";
    tmp(14581) := x"0840";
    tmp(14582) := x"0840";
    tmp(14583) := x"0820";
    tmp(14584) := x"0820";
    tmp(14585) := x"0820";
    tmp(14586) := x"0820";
    tmp(14587) := x"0820";
    tmp(14588) := x"0820";
    tmp(14589) := x"0820";
    tmp(14590) := x"0820";
    tmp(14591) := x"0820";
    tmp(14592) := x"0820";
    tmp(14593) := x"0820";
    tmp(14594) := x"0820";
    tmp(14595) := x"0820";
    tmp(14596) := x"0820";
    tmp(14597) := x"0000";
    tmp(14598) := x"0000";
    tmp(14599) := x"0000";
    tmp(14600) := x"0000";
    tmp(14601) := x"0000";
    tmp(14602) := x"0000";
    tmp(14603) := x"0000";
    tmp(14604) := x"0000";
    tmp(14605) := x"0000";
    tmp(14606) := x"0000";
    tmp(14607) := x"0000";
    tmp(14608) := x"0000";
    tmp(14609) := x"0000";
    tmp(14610) := x"0000";
    tmp(14611) := x"0000";
    tmp(14612) := x"0000";
    tmp(14613) := x"0000";
    tmp(14614) := x"0000";
    tmp(14615) := x"0000";
    tmp(14616) := x"0000";
    tmp(14617) := x"0000";
    tmp(14618) := x"0000";
    tmp(14619) := x"0000";
    tmp(14620) := x"0000";
    tmp(14621) := x"0000";
    tmp(14622) := x"0000";
    tmp(14623) := x"0000";
    tmp(14624) := x"0000";
    tmp(14625) := x"0000";
    tmp(14626) := x"0000";
    tmp(14627) := x"0000";
    tmp(14628) := x"0000";
    tmp(14629) := x"0000";
    tmp(14630) := x"0000";
    tmp(14631) := x"0000";
    tmp(14632) := x"0000";
    tmp(14633) := x"0000";
    tmp(14634) := x"0000";
    tmp(14635) := x"0000";
    tmp(14636) := x"0000";
    tmp(14637) := x"0020";
    tmp(14638) := x"0020";
    tmp(14639) := x"0020";
    tmp(14640) := x"1040";
    tmp(14641) := x"c300";
    tmp(14642) := x"c320";
    tmp(14643) := x"c300";
    tmp(14644) := x"c2e0";
    tmp(14645) := x"c320";
    tmp(14646) := x"cb40";
    tmp(14647) := x"cb40";
    tmp(14648) := x"d360";
    tmp(14649) := x"cb60";
    tmp(14650) := x"cb80";
    tmp(14651) := x"cba0";
    tmp(14652) := x"cb80";
    tmp(14653) := x"d3a0";
    tmp(14654) := x"cba0";
    tmp(14655) := x"d3a0";
    tmp(14656) := x"cb80";
    tmp(14657) := x"cb60";
    tmp(14658) := x"cb40";
    tmp(14659) := x"c300";
    tmp(14660) := x"c2c0";
    tmp(14661) := x"bac0";
    tmp(14662) := x"bac0";
    tmp(14663) := x"b280";
    tmp(14664) := x"a260";
    tmp(14665) := x"9a60";
    tmp(14666) := x"9240";
    tmp(14667) := x"9a60";
    tmp(14668) := x"9a60";
    tmp(14669) := x"9a60";
    tmp(14670) := x"a260";
    tmp(14671) := x"a280";
    tmp(14672) := x"bae0";
    tmp(14673) := x"cb60";
    tmp(14674) := x"c341";
    tmp(14675) := x"c341";
    tmp(14676) := x"b2e0";
    tmp(14677) := x"a260";
    tmp(14678) := x"9a40";
    tmp(14679) := x"9240";
    tmp(14680) := x"a280";
    tmp(14681) := x"a280";
    tmp(14682) := x"aac0";
    tmp(14683) := x"aac0";
    tmp(14684) := x"aac0";
    tmp(14685) := x"a280";
    tmp(14686) := x"a260";
    tmp(14687) := x"aa80";
    tmp(14688) := x"aa80";
    tmp(14689) := x"9a40";
    tmp(14690) := x"9a40";
    tmp(14691) := x"9a40";
    tmp(14692) := x"a260";
    tmp(14693) := x"aa80";
    tmp(14694) := x"a260";
    tmp(14695) := x"aa60";
    tmp(14696) := x"aa80";
    tmp(14697) := x"a260";
    tmp(14698) := x"9220";
    tmp(14699) := x"9220";
    tmp(14700) := x"9200";
    tmp(14701) := x"89e0";
    tmp(14702) := x"7980";
    tmp(14703) := x"7960";
    tmp(14704) := x"7160";
    tmp(14705) := x"7160";
    tmp(14706) := x"6980";
    tmp(14707) := x"7180";
    tmp(14708) := x"79c0";
    tmp(14709) := x"8220";
    tmp(14710) := x"7a00";
    tmp(14711) := x"3920";
    tmp(14712) := x"1080";
    tmp(14713) := x"0860";
    tmp(14714) := x"0840";
    tmp(14715) := x"0840";
    tmp(14716) := x"0020";
    tmp(14717) := x"0000";
    tmp(14718) := x"0000";
    tmp(14719) := x"0000";
    tmp(14720) := x"0000";
    tmp(14721) := x"0000";
    tmp(14722) := x"0000";
    tmp(14723) := x"0000";
    tmp(14724) := x"0000";
    tmp(14725) := x"0000";
    tmp(14726) := x"0000";
    tmp(14727) := x"0000";
    tmp(14728) := x"0000";
    tmp(14729) := x"0000";
    tmp(14730) := x"0000";
    tmp(14731) := x"0000";
    tmp(14732) := x"0000";
    tmp(14733) := x"0000";
    tmp(14734) := x"0000";
    tmp(14735) := x"0000";
    tmp(14736) := x"0000";
    tmp(14737) := x"3964";
    tmp(14738) := x"72ed";
    tmp(14739) := x"6acd";
    tmp(14740) := x"72ad";
    tmp(14741) := x"72ce";
    tmp(14742) := x"7aef";
    tmp(14743) := x"72ad";
    tmp(14744) := x"7aee";
    tmp(14745) := x"9391";
    tmp(14746) := x"9bd3";
    tmp(14747) := x"a455";
    tmp(14748) := x"ac33";
    tmp(14749) := x"ccf7";
    tmp(14750) := x"ee1b";
    tmp(14751) := x"fe9e";
    tmp(14752) := x"edfc";
    tmp(14753) := x"e59b";
    tmp(14754) := x"fe7d";
    tmp(14755) := x"ee1d";
    tmp(14756) := x"ccf9";
    tmp(14757) := x"d579";
    tmp(14758) := x"c454";
    tmp(14759) := x"ee1a";
    tmp(14760) := x"ffdf";
    tmp(14761) := x"eedb";
    tmp(14762) := x"49e7";
    tmp(14763) := x"0020";
    tmp(14764) := x"0000";
    tmp(14765) := x"18a2";
    tmp(14766) := x"ac71";
    tmp(14767) := x"3986";
    tmp(14768) := x"0000";
    tmp(14769) := x"3104";
    tmp(14770) := x"c4d4";
    tmp(14771) := x"6249";
    tmp(14772) := x"0820";
    tmp(14773) := x"8b4d";
    tmp(14774) := x"6aab";
    tmp(14775) := x"1041";
    tmp(14776) := x"a411";
    tmp(14777) := x"6a8a";
    tmp(14778) := x"4165";
    tmp(14779) := x"3945";
    tmp(14780) := x"28a3";
    tmp(14781) := x"3124";
    tmp(14782) := x"82ec";
    tmp(14783) := x"ff9e";
    tmp(14784) := x"736a";
    tmp(14785) := x"10a0";
    tmp(14786) := x"08a0";
    tmp(14787) := x"08a0";
    tmp(14788) := x"08a0";
    tmp(14789) := x"10c0";
    tmp(14790) := x"10c0";
    tmp(14791) := x"1100";
    tmp(14792) := x"1120";
    tmp(14793) := x"1940";
    tmp(14794) := x"2180";
    tmp(14795) := x"2160";
    tmp(14796) := x"21c0";
    tmp(14797) := x"2200";
    tmp(14798) := x"0920";
    tmp(14799) := x"08a0";
    tmp(14800) := x"08c0";
    tmp(14801) := x"08c0";
    tmp(14802) := x"08a0";
    tmp(14803) := x"08c0";
    tmp(14804) := x"08a0";
    tmp(14805) := x"08c0";
    tmp(14806) := x"08a0";
    tmp(14807) := x"08a0";
    tmp(14808) := x"08a0";
    tmp(14809) := x"08a0";
    tmp(14810) := x"08a0";
    tmp(14811) := x"0880";
    tmp(14812) := x"0880";
    tmp(14813) := x"0880";
    tmp(14814) := x"0860";
    tmp(14815) := x"0860";
    tmp(14816) := x"0860";
    tmp(14817) := x"0860";
    tmp(14818) := x"0840";
    tmp(14819) := x"0840";
    tmp(14820) := x"0840";
    tmp(14821) := x"0840";
    tmp(14822) := x"0840";
    tmp(14823) := x"0840";
    tmp(14824) := x"0840";
    tmp(14825) := x"0840";
    tmp(14826) := x"0820";
    tmp(14827) := x"0840";
    tmp(14828) := x"0820";
    tmp(14829) := x"0820";
    tmp(14830) := x"0820";
    tmp(14831) := x"0820";
    tmp(14832) := x"0820";
    tmp(14833) := x"0820";
    tmp(14834) := x"0820";
    tmp(14835) := x"0820";
    tmp(14836) := x"0820";
    tmp(14837) := x"0000";
    tmp(14838) := x"0000";
    tmp(14839) := x"0000";
    tmp(14840) := x"0000";
    tmp(14841) := x"0000";
    tmp(14842) := x"0000";
    tmp(14843) := x"0000";
    tmp(14844) := x"0000";
    tmp(14845) := x"0000";
    tmp(14846) := x"0000";
    tmp(14847) := x"0000";
    tmp(14848) := x"0000";
    tmp(14849) := x"0000";
    tmp(14850) := x"0000";
    tmp(14851) := x"0000";
    tmp(14852) := x"0000";
    tmp(14853) := x"0000";
    tmp(14854) := x"0000";
    tmp(14855) := x"0000";
    tmp(14856) := x"0000";
    tmp(14857) := x"0000";
    tmp(14858) := x"0000";
    tmp(14859) := x"0000";
    tmp(14860) := x"0000";
    tmp(14861) := x"0000";
    tmp(14862) := x"0000";
    tmp(14863) := x"0000";
    tmp(14864) := x"0000";
    tmp(14865) := x"0000";
    tmp(14866) := x"0000";
    tmp(14867) := x"0000";
    tmp(14868) := x"0000";
    tmp(14869) := x"0000";
    tmp(14870) := x"0000";
    tmp(14871) := x"0000";
    tmp(14872) := x"0000";
    tmp(14873) := x"0000";
    tmp(14874) := x"0000";
    tmp(14875) := x"0000";
    tmp(14876) := x"0000";
    tmp(14877) := x"0020";
    tmp(14878) := x"0020";
    tmp(14879) := x"0020";
    tmp(14880) := x"1040";
    tmp(14881) := x"c2e0";
    tmp(14882) := x"c2e0";
    tmp(14883) := x"c2e0";
    tmp(14884) := x"bac0";
    tmp(14885) := x"cb20";
    tmp(14886) := x"cb40";
    tmp(14887) := x"d380";
    tmp(14888) := x"db80";
    tmp(14889) := x"d380";
    tmp(14890) := x"dba0";
    tmp(14891) := x"dbc0";
    tmp(14892) := x"dbc0";
    tmp(14893) := x"dc00";
    tmp(14894) := x"dc00";
    tmp(14895) := x"e3e0";
    tmp(14896) := x"dbe0";
    tmp(14897) := x"d3c0";
    tmp(14898) := x"dba0";
    tmp(14899) := x"db60";
    tmp(14900) := x"d340";
    tmp(14901) := x"cb40";
    tmp(14902) := x"c320";
    tmp(14903) := x"bae0";
    tmp(14904) := x"b2c0";
    tmp(14905) := x"aa80";
    tmp(14906) := x"a280";
    tmp(14907) := x"aaa0";
    tmp(14908) := x"aaa0";
    tmp(14909) := x"aa80";
    tmp(14910) := x"b2c0";
    tmp(14911) := x"aaa0";
    tmp(14912) := x"b2c0";
    tmp(14913) := x"cb40";
    tmp(14914) := x"dba0";
    tmp(14915) := x"d3a1";
    tmp(14916) := x"cb81";
    tmp(14917) := x"b2e0";
    tmp(14918) := x"9a60";
    tmp(14919) := x"9a60";
    tmp(14920) := x"9a60";
    tmp(14921) := x"9a80";
    tmp(14922) := x"9a80";
    tmp(14923) := x"9a80";
    tmp(14924) := x"9a60";
    tmp(14925) := x"9a60";
    tmp(14926) := x"a260";
    tmp(14927) := x"a260";
    tmp(14928) := x"a260";
    tmp(14929) := x"a240";
    tmp(14930) := x"9a40";
    tmp(14931) := x"9a20";
    tmp(14932) := x"9a20";
    tmp(14933) := x"9a20";
    tmp(14934) := x"9a40";
    tmp(14935) := x"a260";
    tmp(14936) := x"a260";
    tmp(14937) := x"9a40";
    tmp(14938) := x"9220";
    tmp(14939) := x"9a20";
    tmp(14940) := x"9200";
    tmp(14941) := x"9200";
    tmp(14942) := x"89c0";
    tmp(14943) := x"89c0";
    tmp(14944) := x"7980";
    tmp(14945) := x"7160";
    tmp(14946) := x"6960";
    tmp(14947) := x"6140";
    tmp(14948) := x"5120";
    tmp(14949) := x"4900";
    tmp(14950) := x"3900";
    tmp(14951) := x"18a0";
    tmp(14952) := x"0860";
    tmp(14953) := x"0840";
    tmp(14954) := x"0840";
    tmp(14955) := x"0020";
    tmp(14956) := x"0020";
    tmp(14957) := x"0000";
    tmp(14958) := x"0000";
    tmp(14959) := x"0000";
    tmp(14960) := x"0000";
    tmp(14961) := x"0000";
    tmp(14962) := x"0000";
    tmp(14963) := x"0000";
    tmp(14964) := x"0000";
    tmp(14965) := x"0000";
    tmp(14966) := x"0000";
    tmp(14967) := x"0000";
    tmp(14968) := x"0000";
    tmp(14969) := x"0000";
    tmp(14970) := x"0000";
    tmp(14971) := x"0000";
    tmp(14972) := x"0000";
    tmp(14973) := x"0000";
    tmp(14974) := x"0000";
    tmp(14975) := x"0000";
    tmp(14976) := x"0820";
    tmp(14977) := x"5a28";
    tmp(14978) := x"624a";
    tmp(14979) := x"6aad";
    tmp(14980) := x"72cd";
    tmp(14981) := x"6aad";
    tmp(14982) := x"6a8c";
    tmp(14983) := x"8b2f";
    tmp(14984) := x"832e";
    tmp(14985) := x"8b50";
    tmp(14986) := x"a3f4";
    tmp(14987) := x"a3d2";
    tmp(14988) := x"cd17";
    tmp(14989) := x"dd59";
    tmp(14990) := x"dd7a";
    tmp(14991) := x"edfc";
    tmp(14992) := x"ee1b";
    tmp(14993) := x"f69d";
    tmp(14994) := x"f67d";
    tmp(14995) := x"e5bb";
    tmp(14996) := x"edbb";
    tmp(14997) := x"d558";
    tmp(14998) := x"dd37";
    tmp(14999) := x"fede";
    tmp(15000) := x"ff1e";
    tmp(15001) := x"eedc";
    tmp(15002) := x"2924";
    tmp(15003) := x"0020";
    tmp(15004) := x"0820";
    tmp(15005) := x"41a6";
    tmp(15006) := x"6acb";
    tmp(15007) := x"0820";
    tmp(15008) := x"1061";
    tmp(15009) := x"938d";
    tmp(15010) := x"c4d4";
    tmp(15011) := x"1041";
    tmp(15012) := x"1881";
    tmp(15013) := x"8b4d";
    tmp(15014) := x"938f";
    tmp(15015) := x"28e3";
    tmp(15016) := x"49c7";
    tmp(15017) := x"28e4";
    tmp(15018) := x"3104";
    tmp(15019) := x"a3cf";
    tmp(15020) := x"728a";
    tmp(15021) := x"20a2";
    tmp(15022) := x"2903";
    tmp(15023) := x"8bad";
    tmp(15024) := x"39a3";
    tmp(15025) := x"08a0";
    tmp(15026) := x"0880";
    tmp(15027) := x"0880";
    tmp(15028) := x"08a0";
    tmp(15029) := x"10c0";
    tmp(15030) := x"10e0";
    tmp(15031) := x"1100";
    tmp(15032) := x"1120";
    tmp(15033) := x"2180";
    tmp(15034) := x"21a0";
    tmp(15035) := x"21a0";
    tmp(15036) := x"2a00";
    tmp(15037) := x"2a60";
    tmp(15038) := x"1120";
    tmp(15039) := x"08a0";
    tmp(15040) := x"08c0";
    tmp(15041) := x"08c0";
    tmp(15042) := x"08c0";
    tmp(15043) := x"08c0";
    tmp(15044) := x"08c0";
    tmp(15045) := x"08c0";
    tmp(15046) := x"08a0";
    tmp(15047) := x"08a0";
    tmp(15048) := x"08c0";
    tmp(15049) := x"08a0";
    tmp(15050) := x"08a0";
    tmp(15051) := x"08a0";
    tmp(15052) := x"08a0";
    tmp(15053) := x"0880";
    tmp(15054) := x"0880";
    tmp(15055) := x"0880";
    tmp(15056) := x"0880";
    tmp(15057) := x"0860";
    tmp(15058) := x"0860";
    tmp(15059) := x"0860";
    tmp(15060) := x"0840";
    tmp(15061) := x"0840";
    tmp(15062) := x"0840";
    tmp(15063) := x"0840";
    tmp(15064) := x"0840";
    tmp(15065) := x"0840";
    tmp(15066) := x"0840";
    tmp(15067) := x"0840";
    tmp(15068) := x"0840";
    tmp(15069) := x"0820";
    tmp(15070) := x"0820";
    tmp(15071) := x"0820";
    tmp(15072) := x"0820";
    tmp(15073) := x"0820";
    tmp(15074) := x"0820";
    tmp(15075) := x"0820";
    tmp(15076) := x"0820";
    tmp(15077) := x"0000";
    tmp(15078) := x"0000";
    tmp(15079) := x"0000";
    tmp(15080) := x"0000";
    tmp(15081) := x"0000";
    tmp(15082) := x"0000";
    tmp(15083) := x"0000";
    tmp(15084) := x"0000";
    tmp(15085) := x"0000";
    tmp(15086) := x"0000";
    tmp(15087) := x"0000";
    tmp(15088) := x"0000";
    tmp(15089) := x"0000";
    tmp(15090) := x"0000";
    tmp(15091) := x"0000";
    tmp(15092) := x"0000";
    tmp(15093) := x"0000";
    tmp(15094) := x"0000";
    tmp(15095) := x"0000";
    tmp(15096) := x"0000";
    tmp(15097) := x"0000";
    tmp(15098) := x"0000";
    tmp(15099) := x"0000";
    tmp(15100) := x"0000";
    tmp(15101) := x"0000";
    tmp(15102) := x"0000";
    tmp(15103) := x"0000";
    tmp(15104) := x"0000";
    tmp(15105) := x"0000";
    tmp(15106) := x"0000";
    tmp(15107) := x"0000";
    tmp(15108) := x"0000";
    tmp(15109) := x"0000";
    tmp(15110) := x"0000";
    tmp(15111) := x"0000";
    tmp(15112) := x"0000";
    tmp(15113) := x"0000";
    tmp(15114) := x"0000";
    tmp(15115) := x"0000";
    tmp(15116) := x"0000";
    tmp(15117) := x"0020";
    tmp(15118) := x"0020";
    tmp(15119) := x"0020";
    tmp(15120) := x"1040";
    tmp(15121) := x"c2c0";
    tmp(15122) := x"bac0";
    tmp(15123) := x"bac0";
    tmp(15124) := x"c2e0";
    tmp(15125) := x"cb20";
    tmp(15126) := x"cb40";
    tmp(15127) := x"db80";
    tmp(15128) := x"db80";
    tmp(15129) := x"dba0";
    tmp(15130) := x"dba0";
    tmp(15131) := x"e3c0";
    tmp(15132) := x"d380";
    tmp(15133) := x"d3a0";
    tmp(15134) := x"cb80";
    tmp(15135) := x"d380";
    tmp(15136) := x"cb40";
    tmp(15137) := x"c340";
    tmp(15138) := x"cb20";
    tmp(15139) := x"cb20";
    tmp(15140) := x"cb20";
    tmp(15141) := x"d340";
    tmp(15142) := x"cb40";
    tmp(15143) := x"c320";
    tmp(15144) := x"c300";
    tmp(15145) := x"bac0";
    tmp(15146) := x"b2c0";
    tmp(15147) := x"b2c0";
    tmp(15148) := x"bae0";
    tmp(15149) := x"bac0";
    tmp(15150) := x"bae0";
    tmp(15151) := x"bac0";
    tmp(15152) := x"bac0";
    tmp(15153) := x"bae0";
    tmp(15154) := x"c320";
    tmp(15155) := x"cb80";
    tmp(15156) := x"dbe0";
    tmp(15157) := x"cb60";
    tmp(15158) := x"aac0";
    tmp(15159) := x"9a60";
    tmp(15160) := x"9a60";
    tmp(15161) := x"9a60";
    tmp(15162) := x"9a60";
    tmp(15163) := x"9a60";
    tmp(15164) := x"9a80";
    tmp(15165) := x"9a60";
    tmp(15166) := x"a260";
    tmp(15167) := x"a260";
    tmp(15168) := x"a240";
    tmp(15169) := x"a260";
    tmp(15170) := x"a240";
    tmp(15171) := x"a240";
    tmp(15172) := x"a240";
    tmp(15173) := x"9a40";
    tmp(15174) := x"9a20";
    tmp(15175) := x"9220";
    tmp(15176) := x"9220";
    tmp(15177) := x"9a20";
    tmp(15178) := x"9a20";
    tmp(15179) := x"a220";
    tmp(15180) := x"9a20";
    tmp(15181) := x"9200";
    tmp(15182) := x"9200";
    tmp(15183) := x"89e0";
    tmp(15184) := x"81c0";
    tmp(15185) := x"7180";
    tmp(15186) := x"6960";
    tmp(15187) := x"5920";
    tmp(15188) := x"4900";
    tmp(15189) := x"38e0";
    tmp(15190) := x"20a0";
    tmp(15191) := x"1080";
    tmp(15192) := x"0840";
    tmp(15193) := x"0840";
    tmp(15194) := x"0020";
    tmp(15195) := x"0020";
    tmp(15196) := x"0020";
    tmp(15197) := x"0000";
    tmp(15198) := x"0000";
    tmp(15199) := x"0000";
    tmp(15200) := x"0000";
    tmp(15201) := x"0000";
    tmp(15202) := x"0000";
    tmp(15203) := x"0000";
    tmp(15204) := x"0000";
    tmp(15205) := x"0000";
    tmp(15206) := x"0000";
    tmp(15207) := x"0000";
    tmp(15208) := x"0000";
    tmp(15209) := x"0000";
    tmp(15210) := x"0000";
    tmp(15211) := x"0000";
    tmp(15212) := x"0000";
    tmp(15213) := x"0000";
    tmp(15214) := x"0000";
    tmp(15215) := x"0000";
    tmp(15216) := x"20a2";
    tmp(15217) := x"5a08";
    tmp(15218) := x"5a29";
    tmp(15219) := x"728d";
    tmp(15220) := x"728c";
    tmp(15221) := x"7acd";
    tmp(15222) := x"7acd";
    tmp(15223) := x"7aad";
    tmp(15224) := x"93b1";
    tmp(15225) := x"8b0f";
    tmp(15226) := x"934f";
    tmp(15227) := x"bc32";
    tmp(15228) := x"ccd6";
    tmp(15229) := x"c496";
    tmp(15230) := x"dd39";
    tmp(15231) := x"edfd";
    tmp(15232) := x"ee7d";
    tmp(15233) := x"ee3c";
    tmp(15234) := x"edfb";
    tmp(15235) := x"edfb";
    tmp(15236) := x"fe3d";
    tmp(15237) := x"dd38";
    tmp(15238) := x"f6bc";
    tmp(15239) := x"fedd";
    tmp(15240) := x"e579";
    tmp(15241) := x"5a4a";
    tmp(15242) := x"0841";
    tmp(15243) := x"0820";
    tmp(15244) := x"3144";
    tmp(15245) := x"9c51";
    tmp(15246) := x"1882";
    tmp(15247) := x"0020";
    tmp(15248) := x"6248";
    tmp(15249) := x"9baf";
    tmp(15250) := x"28c3";
    tmp(15251) := x"0820";
    tmp(15252) := x"6aaa";
    tmp(15253) := x"3125";
    tmp(15254) := x"936f";
    tmp(15255) := x"8b8d";
    tmp(15256) := x"1882";
    tmp(15257) := x"20c3";
    tmp(15258) := x"1882";
    tmp(15259) := x"1882";
    tmp(15260) := x"6249";
    tmp(15261) := x"b491";
    tmp(15262) := x"2903";
    tmp(15263) := x"18a2";
    tmp(15264) := x"10a1";
    tmp(15265) := x"0880";
    tmp(15266) := x"08a0";
    tmp(15267) := x"08a0";
    tmp(15268) := x"0880";
    tmp(15269) := x"10c0";
    tmp(15270) := x"10e0";
    tmp(15271) := x"1100";
    tmp(15272) := x"1920";
    tmp(15273) := x"2180";
    tmp(15274) := x"2180";
    tmp(15275) := x"21a0";
    tmp(15276) := x"2a00";
    tmp(15277) := x"2a20";
    tmp(15278) := x"08e0";
    tmp(15279) := x"08a0";
    tmp(15280) := x"08a0";
    tmp(15281) := x"08a0";
    tmp(15282) := x"08c0";
    tmp(15283) := x"08c0";
    tmp(15284) := x"08c0";
    tmp(15285) := x"08c0";
    tmp(15286) := x"08c0";
    tmp(15287) := x"08c0";
    tmp(15288) := x"08c0";
    tmp(15289) := x"08c0";
    tmp(15290) := x"08c0";
    tmp(15291) := x"08a0";
    tmp(15292) := x"08a0";
    tmp(15293) := x"08a0";
    tmp(15294) := x"08a0";
    tmp(15295) := x"0880";
    tmp(15296) := x"0880";
    tmp(15297) := x"0880";
    tmp(15298) := x"0860";
    tmp(15299) := x"0860";
    tmp(15300) := x"0860";
    tmp(15301) := x"0860";
    tmp(15302) := x"0860";
    tmp(15303) := x"0840";
    tmp(15304) := x"0840";
    tmp(15305) := x"0840";
    tmp(15306) := x"0840";
    tmp(15307) := x"0840";
    tmp(15308) := x"0840";
    tmp(15309) := x"0840";
    tmp(15310) := x"0840";
    tmp(15311) := x"0820";
    tmp(15312) := x"0820";
    tmp(15313) := x"0820";
    tmp(15314) := x"0820";
    tmp(15315) := x"0820";
    tmp(15316) := x"0820";
    tmp(15317) := x"0000";
    tmp(15318) := x"0000";
    tmp(15319) := x"0000";
    tmp(15320) := x"0000";
    tmp(15321) := x"0000";
    tmp(15322) := x"0000";
    tmp(15323) := x"0000";
    tmp(15324) := x"0000";
    tmp(15325) := x"0000";
    tmp(15326) := x"0000";
    tmp(15327) := x"0000";
    tmp(15328) := x"0000";
    tmp(15329) := x"0000";
    tmp(15330) := x"0000";
    tmp(15331) := x"0000";
    tmp(15332) := x"0000";
    tmp(15333) := x"0000";
    tmp(15334) := x"0000";
    tmp(15335) := x"0000";
    tmp(15336) := x"0000";
    tmp(15337) := x"0000";
    tmp(15338) := x"0000";
    tmp(15339) := x"0000";
    tmp(15340) := x"0000";
    tmp(15341) := x"0000";
    tmp(15342) := x"0000";
    tmp(15343) := x"0000";
    tmp(15344) := x"0000";
    tmp(15345) := x"0000";
    tmp(15346) := x"0000";
    tmp(15347) := x"0000";
    tmp(15348) := x"0000";
    tmp(15349) := x"0000";
    tmp(15350) := x"0000";
    tmp(15351) := x"0000";
    tmp(15352) := x"0000";
    tmp(15353) := x"0000";
    tmp(15354) := x"0000";
    tmp(15355) := x"0000";
    tmp(15356) := x"0000";
    tmp(15357) := x"0020";
    tmp(15358) := x"0020";
    tmp(15359) := x"0020";
    tmp(15360) := x"1040";
    tmp(15361) := x"bac0";
    tmp(15362) := x"bac0";
    tmp(15363) := x"bae0";
    tmp(15364) := x"c300";
    tmp(15365) := x"c320";
    tmp(15366) := x"cb40";
    tmp(15367) := x"cb40";
    tmp(15368) := x"cb20";
    tmp(15369) := x"c300";
    tmp(15370) := x"cb40";
    tmp(15371) := x"cb40";
    tmp(15372) := x"cb20";
    tmp(15373) := x"cb20";
    tmp(15374) := x"bb00";
    tmp(15375) := x"bae0";
    tmp(15376) := x"c300";
    tmp(15377) := x"c300";
    tmp(15378) := x"cb20";
    tmp(15379) := x"c320";
    tmp(15380) := x"cb00";
    tmp(15381) := x"cb00";
    tmp(15382) := x"cb00";
    tmp(15383) := x"c2e0";
    tmp(15384) := x"cae0";
    tmp(15385) := x"c2e0";
    tmp(15386) := x"c2e0";
    tmp(15387) := x"cb20";
    tmp(15388) := x"d340";
    tmp(15389) := x"d340";
    tmp(15390) := x"cb20";
    tmp(15391) := x"cb40";
    tmp(15392) := x"d340";
    tmp(15393) := x"d360";
    tmp(15394) := x"cb40";
    tmp(15395) := x"d380";
    tmp(15396) := x"dbc0";
    tmp(15397) := x"cb60";
    tmp(15398) := x"b2c0";
    tmp(15399) := x"9a80";
    tmp(15400) := x"a280";
    tmp(15401) := x"a280";
    tmp(15402) := x"a260";
    tmp(15403) := x"a260";
    tmp(15404) := x"a2a0";
    tmp(15405) := x"aaa0";
    tmp(15406) := x"aa80";
    tmp(15407) := x"9a60";
    tmp(15408) := x"a240";
    tmp(15409) := x"9a20";
    tmp(15410) := x"a220";
    tmp(15411) := x"9a40";
    tmp(15412) := x"9a40";
    tmp(15413) := x"9a20";
    tmp(15414) := x"9a20";
    tmp(15415) := x"9a20";
    tmp(15416) := x"9a40";
    tmp(15417) := x"9a40";
    tmp(15418) := x"a240";
    tmp(15419) := x"a240";
    tmp(15420) := x"a260";
    tmp(15421) := x"a220";
    tmp(15422) := x"9a20";
    tmp(15423) := x"9200";
    tmp(15424) := x"89c0";
    tmp(15425) := x"79a0";
    tmp(15426) := x"6980";
    tmp(15427) := x"6140";
    tmp(15428) := x"5120";
    tmp(15429) := x"30e0";
    tmp(15430) := x"1880";
    tmp(15431) := x"0860";
    tmp(15432) := x"0840";
    tmp(15433) := x"0020";
    tmp(15434) := x"0020";
    tmp(15435) := x"0020";
    tmp(15436) := x"0020";
    tmp(15437) := x"0020";
    tmp(15438) := x"0020";
    tmp(15439) := x"0000";
    tmp(15440) := x"0000";
    tmp(15441) := x"0000";
    tmp(15442) := x"0000";
    tmp(15443) := x"0000";
    tmp(15444) := x"0000";
    tmp(15445) := x"0000";
    tmp(15446) := x"0000";
    tmp(15447) := x"0000";
    tmp(15448) := x"0000";
    tmp(15449) := x"0000";
    tmp(15450) := x"0000";
    tmp(15451) := x"0000";
    tmp(15452) := x"0000";
    tmp(15453) := x"0000";
    tmp(15454) := x"0000";
    tmp(15455) := x"0840";
    tmp(15456) := x"5a27";
    tmp(15457) := x"51e7";
    tmp(15458) := x"5a09";
    tmp(15459) := x"728c";
    tmp(15460) := x"6a4a";
    tmp(15461) := x"8aee";
    tmp(15462) := x"8b0e";
    tmp(15463) := x"82ee";
    tmp(15464) := x"7acd";
    tmp(15465) := x"930e";
    tmp(15466) := x"abd1";
    tmp(15467) := x"bc54";
    tmp(15468) := x"b413";
    tmp(15469) := x"c496";
    tmp(15470) := x"dd39";
    tmp(15471) := x"edfb";
    tmp(15472) := x"f69e";
    tmp(15473) := x"ee3c";
    tmp(15474) := x"ee9d";
    tmp(15475) := x"ee5c";
    tmp(15476) := x"edba";
    tmp(15477) := x"ed99";
    tmp(15478) := x"ff7e";
    tmp(15479) := x"e578";
    tmp(15480) := x"ed98";
    tmp(15481) := x"3966";
    tmp(15482) := x"0020";
    tmp(15483) := x"18a2";
    tmp(15484) := x"9bf0";
    tmp(15485) := x"4a07";
    tmp(15486) := x"0000";
    tmp(15487) := x"28e3";
    tmp(15488) := x"d555";
    tmp(15489) := x"20c3";
    tmp(15490) := x"0820";
    tmp(15491) := x"2903";
    tmp(15492) := x"938f";
    tmp(15493) := x"20a3";
    tmp(15494) := x"834e";
    tmp(15495) := x"1882";
    tmp(15496) := x"5208";
    tmp(15497) := x"3966";
    tmp(15498) := x"8b8e";
    tmp(15499) := x"3125";
    tmp(15500) := x"1882";
    tmp(15501) := x"20a2";
    tmp(15502) := x"5207";
    tmp(15503) := x"18a1";
    tmp(15504) := x"0840";
    tmp(15505) := x"0860";
    tmp(15506) := x"08a0";
    tmp(15507) := x"08c0";
    tmp(15508) := x"10c0";
    tmp(15509) := x"10e0";
    tmp(15510) := x"1100";
    tmp(15511) := x"1920";
    tmp(15512) := x"1920";
    tmp(15513) := x"21a0";
    tmp(15514) := x"21a0";
    tmp(15515) := x"21c0";
    tmp(15516) := x"2200";
    tmp(15517) := x"19a0";
    tmp(15518) := x"08a0";
    tmp(15519) := x"08a0";
    tmp(15520) := x"08a0";
    tmp(15521) := x"08a0";
    tmp(15522) := x"08a0";
    tmp(15523) := x"08a0";
    tmp(15524) := x"08c0";
    tmp(15525) := x"08c0";
    tmp(15526) := x"08c0";
    tmp(15527) := x"08c0";
    tmp(15528) := x"08c0";
    tmp(15529) := x"08c0";
    tmp(15530) := x"08c0";
    tmp(15531) := x"08c0";
    tmp(15532) := x"08a0";
    tmp(15533) := x"08a0";
    tmp(15534) := x"08a0";
    tmp(15535) := x"08a0";
    tmp(15536) := x"08a0";
    tmp(15537) := x"0880";
    tmp(15538) := x"0880";
    tmp(15539) := x"0880";
    tmp(15540) := x"0860";
    tmp(15541) := x"0860";
    tmp(15542) := x"0860";
    tmp(15543) := x"0860";
    tmp(15544) := x"0860";
    tmp(15545) := x"0840";
    tmp(15546) := x"0840";
    tmp(15547) := x"0840";
    tmp(15548) := x"0840";
    tmp(15549) := x"0840";
    tmp(15550) := x"0840";
    tmp(15551) := x"0840";
    tmp(15552) := x"0820";
    tmp(15553) := x"0820";
    tmp(15554) := x"0820";
    tmp(15555) := x"0820";
    tmp(15556) := x"0820";
    tmp(15557) := x"0000";
    tmp(15558) := x"0000";
    tmp(15559) := x"0000";
    tmp(15560) := x"0000";
    tmp(15561) := x"0000";
    tmp(15562) := x"0000";
    tmp(15563) := x"0000";
    tmp(15564) := x"0000";
    tmp(15565) := x"0000";
    tmp(15566) := x"0000";
    tmp(15567) := x"0000";
    tmp(15568) := x"0000";
    tmp(15569) := x"0000";
    tmp(15570) := x"0000";
    tmp(15571) := x"0000";
    tmp(15572) := x"0000";
    tmp(15573) := x"0000";
    tmp(15574) := x"0000";
    tmp(15575) := x"0000";
    tmp(15576) := x"0000";
    tmp(15577) := x"0000";
    tmp(15578) := x"0000";
    tmp(15579) := x"0000";
    tmp(15580) := x"0000";
    tmp(15581) := x"0000";
    tmp(15582) := x"0000";
    tmp(15583) := x"0000";
    tmp(15584) := x"0000";
    tmp(15585) := x"0000";
    tmp(15586) := x"0000";
    tmp(15587) := x"0000";
    tmp(15588) := x"0000";
    tmp(15589) := x"0000";
    tmp(15590) := x"0000";
    tmp(15591) := x"0000";
    tmp(15592) := x"0000";
    tmp(15593) := x"0000";
    tmp(15594) := x"0000";
    tmp(15595) := x"0000";
    tmp(15596) := x"0000";
    tmp(15597) := x"0020";
    tmp(15598) := x"0020";
    tmp(15599) := x"0020";
    tmp(15600) := x"1040";
    tmp(15601) := x"bac0";
    tmp(15602) := x"b2c0";
    tmp(15603) := x"b2e0";
    tmp(15604) := x"bb00";
    tmp(15605) := x"bae0";
    tmp(15606) := x"bae0";
    tmp(15607) := x"c2e0";
    tmp(15608) := x"bac0";
    tmp(15609) := x"bac0";
    tmp(15610) := x"c2e0";
    tmp(15611) := x"bac0";
    tmp(15612) := x"c2c0";
    tmp(15613) := x"cb00";
    tmp(15614) := x"cb20";
    tmp(15615) := x"c2c0";
    tmp(15616) := x"bac0";
    tmp(15617) := x"cb20";
    tmp(15618) := x"db40";
    tmp(15619) := x"cb20";
    tmp(15620) := x"cb20";
    tmp(15621) := x"d320";
    tmp(15622) := x"d300";
    tmp(15623) := x"d2e0";
    tmp(15624) := x"d320";
    tmp(15625) := x"d320";
    tmp(15626) := x"e360";
    tmp(15627) := x"db60";
    tmp(15628) := x"e360";
    tmp(15629) := x"eba0";
    tmp(15630) := x"e380";
    tmp(15631) := x"e3a0";
    tmp(15632) := x"e380";
    tmp(15633) := x"e3a0";
    tmp(15634) := x"ebc0";
    tmp(15635) := x"ec00";
    tmp(15636) := x"e400";
    tmp(15637) := x"d380";
    tmp(15638) := x"b2c0";
    tmp(15639) := x"9a60";
    tmp(15640) := x"9a40";
    tmp(15641) := x"9a40";
    tmp(15642) := x"9a60";
    tmp(15643) := x"aa80";
    tmp(15644) := x"b2c0";
    tmp(15645) := x"b2c0";
    tmp(15646) := x"a260";
    tmp(15647) := x"9a40";
    tmp(15648) := x"a240";
    tmp(15649) := x"a220";
    tmp(15650) := x"9a20";
    tmp(15651) := x"9a20";
    tmp(15652) := x"9200";
    tmp(15653) := x"91e0";
    tmp(15654) := x"9a20";
    tmp(15655) := x"9a20";
    tmp(15656) := x"9220";
    tmp(15657) := x"a240";
    tmp(15658) := x"aa60";
    tmp(15659) := x"aa60";
    tmp(15660) := x"b280";
    tmp(15661) := x"aa40";
    tmp(15662) := x"a220";
    tmp(15663) := x"91e0";
    tmp(15664) := x"81a0";
    tmp(15665) := x"79a0";
    tmp(15666) := x"6980";
    tmp(15667) := x"5960";
    tmp(15668) := x"4920";
    tmp(15669) := x"28c0";
    tmp(15670) := x"1880";
    tmp(15671) := x"0840";
    tmp(15672) := x"0020";
    tmp(15673) := x"0020";
    tmp(15674) := x"0020";
    tmp(15675) := x"0020";
    tmp(15676) := x"0020";
    tmp(15677) := x"0020";
    tmp(15678) := x"0020";
    tmp(15679) := x"0020";
    tmp(15680) := x"0020";
    tmp(15681) := x"0000";
    tmp(15682) := x"0000";
    tmp(15683) := x"0000";
    tmp(15684) := x"0000";
    tmp(15685) := x"0000";
    tmp(15686) := x"0000";
    tmp(15687) := x"0000";
    tmp(15688) := x"0000";
    tmp(15689) := x"0000";
    tmp(15690) := x"0000";
    tmp(15691) := x"0000";
    tmp(15692) := x"0000";
    tmp(15693) := x"0000";
    tmp(15694) := x"0820";
    tmp(15695) := x"41a5";
    tmp(15696) := x"72cb";
    tmp(15697) := x"6228";
    tmp(15698) := x"7acc";
    tmp(15699) := x"8b2e";
    tmp(15700) := x"728b";
    tmp(15701) := x"7acd";
    tmp(15702) := x"82ee";
    tmp(15703) := x"82ee";
    tmp(15704) := x"8b2e";
    tmp(15705) := x"b412";
    tmp(15706) := x"b433";
    tmp(15707) := x"a3b2";
    tmp(15708) := x"9b71";
    tmp(15709) := x"bc54";
    tmp(15710) := x"ccf7";
    tmp(15711) := x"f65d";
    tmp(15712) := x"ee3d";
    tmp(15713) := x"eedd";
    tmp(15714) := x"ee3c";
    tmp(15715) := x"f65d";
    tmp(15716) := x"f69c";
    tmp(15717) := x"fe9d";
    tmp(15718) := x"ff3e";
    tmp(15719) := x"e516";
    tmp(15720) := x"bcf5";
    tmp(15721) := x"0821";
    tmp(15722) := x"0820";
    tmp(15723) := x"5a49";
    tmp(15724) := x"93f0";
    tmp(15725) := x"0820";
    tmp(15726) := x"0020";
    tmp(15727) := x"6a69";
    tmp(15728) := x"b4b3";
    tmp(15729) := x"0841";
    tmp(15730) := x"28e3";
    tmp(15731) := x"9c10";
    tmp(15732) := x"20a3";
    tmp(15733) := x"28e4";
    tmp(15734) := x"730c";
    tmp(15735) := x"28e4";
    tmp(15736) := x"0821";
    tmp(15737) := x"20c3";
    tmp(15738) := x"936f";
    tmp(15739) := x"bc93";
    tmp(15740) := x"9bcf";
    tmp(15741) := x"3965";
    tmp(15742) := x"1862";
    tmp(15743) := x"3123";
    tmp(15744) := x"10a0";
    tmp(15745) := x"0860";
    tmp(15746) := x"08c0";
    tmp(15747) := x"10e0";
    tmp(15748) := x"10c0";
    tmp(15749) := x"10c0";
    tmp(15750) := x"1100";
    tmp(15751) := x"10e0";
    tmp(15752) := x"1920";
    tmp(15753) := x"21a0";
    tmp(15754) := x"21a0";
    tmp(15755) := x"21e0";
    tmp(15756) := x"2a61";
    tmp(15757) := x"19e1";
    tmp(15758) := x"08a0";
    tmp(15759) := x"08a0";
    tmp(15760) := x"08a0";
    tmp(15761) := x"08a0";
    tmp(15762) := x"08c0";
    tmp(15763) := x"08c0";
    tmp(15764) := x"08c0";
    tmp(15765) := x"08e0";
    tmp(15766) := x"08c0";
    tmp(15767) := x"08e0";
    tmp(15768) := x"08e0";
    tmp(15769) := x"08e0";
    tmp(15770) := x"08e0";
    tmp(15771) := x"08e0";
    tmp(15772) := x"08e0";
    tmp(15773) := x"08c0";
    tmp(15774) := x"08a0";
    tmp(15775) := x"08a0";
    tmp(15776) := x"08a0";
    tmp(15777) := x"08a0";
    tmp(15778) := x"0880";
    tmp(15779) := x"0880";
    tmp(15780) := x"0880";
    tmp(15781) := x"0880";
    tmp(15782) := x"0880";
    tmp(15783) := x"0860";
    tmp(15784) := x"0860";
    tmp(15785) := x"0860";
    tmp(15786) := x"0860";
    tmp(15787) := x"0840";
    tmp(15788) := x"0840";
    tmp(15789) := x"0840";
    tmp(15790) := x"0840";
    tmp(15791) := x"0840";
    tmp(15792) := x"0840";
    tmp(15793) := x"0820";
    tmp(15794) := x"0820";
    tmp(15795) := x"0820";
    tmp(15796) := x"0820";
    tmp(15797) := x"0000";
    tmp(15798) := x"0000";
    tmp(15799) := x"0000";
    tmp(15800) := x"0000";
    tmp(15801) := x"0000";
    tmp(15802) := x"0000";
    tmp(15803) := x"0000";
    tmp(15804) := x"0000";
    tmp(15805) := x"0000";
    tmp(15806) := x"0000";
    tmp(15807) := x"0000";
    tmp(15808) := x"0000";
    tmp(15809) := x"0000";
    tmp(15810) := x"0000";
    tmp(15811) := x"0000";
    tmp(15812) := x"0000";
    tmp(15813) := x"0000";
    tmp(15814) := x"0000";
    tmp(15815) := x"0000";
    tmp(15816) := x"0000";
    tmp(15817) := x"0000";
    tmp(15818) := x"0000";
    tmp(15819) := x"0000";
    tmp(15820) := x"0000";
    tmp(15821) := x"0000";
    tmp(15822) := x"0000";
    tmp(15823) := x"0000";
    tmp(15824) := x"0000";
    tmp(15825) := x"0000";
    tmp(15826) := x"0000";
    tmp(15827) := x"0000";
    tmp(15828) := x"0000";
    tmp(15829) := x"0000";
    tmp(15830) := x"0000";
    tmp(15831) := x"0000";
    tmp(15832) := x"0000";
    tmp(15833) := x"0000";
    tmp(15834) := x"0000";
    tmp(15835) := x"0000";
    tmp(15836) := x"0000";
    tmp(15837) := x"0820";
    tmp(15838) := x"0820";
    tmp(15839) := x"0820";
    tmp(15840) := x"1040";
    tmp(15841) := x"c2e0";
    tmp(15842) := x"b2c0";
    tmp(15843) := x"bae0";
    tmp(15844) := x"b2c0";
    tmp(15845) := x"bac0";
    tmp(15846) := x"bac0";
    tmp(15847) := x"c2e0";
    tmp(15848) := x"baa0";
    tmp(15849) := x"c2c0";
    tmp(15850) := x"c2e0";
    tmp(15851) := x"cb00";
    tmp(15852) := x"cb00";
    tmp(15853) := x"c300";
    tmp(15854) := x"c2c0";
    tmp(15855) := x"c2c0";
    tmp(15856) := x"c2e0";
    tmp(15857) := x"cb20";
    tmp(15858) := x"cb20";
    tmp(15859) := x"d300";
    tmp(15860) := x"d300";
    tmp(15861) := x"d300";
    tmp(15862) := x"d2e0";
    tmp(15863) := x"d2e0";
    tmp(15864) := x"d300";
    tmp(15865) := x"db40";
    tmp(15866) := x"eb60";
    tmp(15867) := x"eb80";
    tmp(15868) := x"eb80";
    tmp(15869) := x"f3c0";
    tmp(15870) := x"f3c0";
    tmp(15871) := x"f3c0";
    tmp(15872) := x"ebc0";
    tmp(15873) := x"f3e0";
    tmp(15874) := x"ebe0";
    tmp(15875) := x"f440";
    tmp(15876) := x"dbc0";
    tmp(15877) := x"bb00";
    tmp(15878) := x"aa80";
    tmp(15879) := x"9a20";
    tmp(15880) := x"9220";
    tmp(15881) := x"9220";
    tmp(15882) := x"aa80";
    tmp(15883) := x"b2c0";
    tmp(15884) := x"bae0";
    tmp(15885) := x"b2c0";
    tmp(15886) := x"aa60";
    tmp(15887) := x"a240";
    tmp(15888) := x"a220";
    tmp(15889) := x"9a00";
    tmp(15890) := x"91e0";
    tmp(15891) := x"9a00";
    tmp(15892) := x"9a00";
    tmp(15893) := x"9200";
    tmp(15894) := x"a220";
    tmp(15895) := x"9a20";
    tmp(15896) := x"9a20";
    tmp(15897) := x"a240";
    tmp(15898) := x"aa60";
    tmp(15899) := x"b280";
    tmp(15900) := x"b280";
    tmp(15901) := x"aa60";
    tmp(15902) := x"a240";
    tmp(15903) := x"91e0";
    tmp(15904) := x"81a0";
    tmp(15905) := x"7180";
    tmp(15906) := x"6980";
    tmp(15907) := x"5140";
    tmp(15908) := x"3100";
    tmp(15909) := x"20c0";
    tmp(15910) := x"1060";
    tmp(15911) := x"0820";
    tmp(15912) := x"0000";
    tmp(15913) := x"0000";
    tmp(15914) := x"0000";
    tmp(15915) := x"0020";
    tmp(15916) := x"0000";
    tmp(15917) := x"0000";
    tmp(15918) := x"0000";
    tmp(15919) := x"0000";
    tmp(15920) := x"0000";
    tmp(15921) := x"0000";
    tmp(15922) := x"0000";
    tmp(15923) := x"0000";
    tmp(15924) := x"0000";
    tmp(15925) := x"0000";
    tmp(15926) := x"0000";
    tmp(15927) := x"0000";
    tmp(15928) := x"0000";
    tmp(15929) := x"0000";
    tmp(15930) := x"0000";
    tmp(15931) := x"0000";
    tmp(15932) := x"0000";
    tmp(15933) := x"0000";
    tmp(15934) := x"20c2";
    tmp(15935) := x"6249";
    tmp(15936) := x"6a8b";
    tmp(15937) := x"82ed";
    tmp(15938) := x"9391";
    tmp(15939) := x"9350";
    tmp(15940) := x"9b90";
    tmp(15941) := x"936f";
    tmp(15942) := x"7a8b";
    tmp(15943) := x"9b70";
    tmp(15944) := x"b433";
    tmp(15945) := x"ac34";
    tmp(15946) := x"9bd2";
    tmp(15947) := x"9370";
    tmp(15948) := x"930f";
    tmp(15949) := x"abd1";
    tmp(15950) := x"dd79";
    tmp(15951) := x"edfc";
    tmp(15952) := x"ee3c";
    tmp(15953) := x"febe";
    tmp(15954) := x"f63c";
    tmp(15955) := x"ff1d";
    tmp(15956) := x"f69c";
    tmp(15957) := x"febc";
    tmp(15958) := x"ff3e";
    tmp(15959) := x"fdd8";
    tmp(15960) := x"3124";
    tmp(15961) := x"0000";
    tmp(15962) := x"0020";
    tmp(15963) := x"938e";
    tmp(15964) := x"5a49";
    tmp(15965) := x"0820";
    tmp(15966) := x"1041";
    tmp(15967) := x"bc92";
    tmp(15968) := x"3965";
    tmp(15969) := x"1061";
    tmp(15970) := x"5a28";
    tmp(15971) := x"d596";
    tmp(15972) := x"0820";
    tmp(15973) := x"4a08";
    tmp(15974) := x"93f1";
    tmp(15975) := x"a492";
    tmp(15976) := x"2904";
    tmp(15977) := x"0820";
    tmp(15978) := x"0821";
    tmp(15979) := x"51e8";
    tmp(15980) := x"832d";
    tmp(15981) := x"49c7";
    tmp(15982) := x"732c";
    tmp(15983) := x"18c2";
    tmp(15984) := x"0840";
    tmp(15985) := x"0880";
    tmp(15986) := x"08a0";
    tmp(15987) := x"10e0";
    tmp(15988) := x"10c0";
    tmp(15989) := x"10c0";
    tmp(15990) := x"10e0";
    tmp(15991) := x"1940";
    tmp(15992) := x"1960";
    tmp(15993) := x"21e0";
    tmp(15994) := x"1980";
    tmp(15995) := x"21e0";
    tmp(15996) := x"32e1";
    tmp(15997) := x"19a1";
    tmp(15998) := x"0880";
    tmp(15999) := x"08a0";
    tmp(16000) := x"08a0";
    tmp(16001) := x"08a0";
    tmp(16002) := x"08c0";
    tmp(16003) := x"08c0";
    tmp(16004) := x"08e0";
    tmp(16005) := x"08e0";
    tmp(16006) := x"08e0";
    tmp(16007) := x"08e0";
    tmp(16008) := x"0900";
    tmp(16009) := x"08e0";
    tmp(16010) := x"0900";
    tmp(16011) := x"0900";
    tmp(16012) := x"08e0";
    tmp(16013) := x"08e0";
    tmp(16014) := x"08e0";
    tmp(16015) := x"08e0";
    tmp(16016) := x"08c0";
    tmp(16017) := x"08a0";
    tmp(16018) := x"08a0";
    tmp(16019) := x"0880";
    tmp(16020) := x"0880";
    tmp(16021) := x"0880";
    tmp(16022) := x"0880";
    tmp(16023) := x"0880";
    tmp(16024) := x"0860";
    tmp(16025) := x"0860";
    tmp(16026) := x"0860";
    tmp(16027) := x"0860";
    tmp(16028) := x"0840";
    tmp(16029) := x"0840";
    tmp(16030) := x"0840";
    tmp(16031) := x"0840";
    tmp(16032) := x"0840";
    tmp(16033) := x"0840";
    tmp(16034) := x"0820";
    tmp(16035) := x"0820";
    tmp(16036) := x"0820";
    tmp(16037) := x"0000";
    tmp(16038) := x"0000";
    tmp(16039) := x"0000";
    tmp(16040) := x"0000";
    tmp(16041) := x"0000";
    tmp(16042) := x"0000";
    tmp(16043) := x"0000";
    tmp(16044) := x"0000";
    tmp(16045) := x"0000";
    tmp(16046) := x"0000";
    tmp(16047) := x"0000";
    tmp(16048) := x"0000";
    tmp(16049) := x"0000";
    tmp(16050) := x"0000";
    tmp(16051) := x"0000";
    tmp(16052) := x"0000";
    tmp(16053) := x"0000";
    tmp(16054) := x"0000";
    tmp(16055) := x"0000";
    tmp(16056) := x"0000";
    tmp(16057) := x"0000";
    tmp(16058) := x"0000";
    tmp(16059) := x"0000";
    tmp(16060) := x"0000";
    tmp(16061) := x"0000";
    tmp(16062) := x"0000";
    tmp(16063) := x"0000";
    tmp(16064) := x"0000";
    tmp(16065) := x"0000";
    tmp(16066) := x"0000";
    tmp(16067) := x"0000";
    tmp(16068) := x"0000";
    tmp(16069) := x"0000";
    tmp(16070) := x"0000";
    tmp(16071) := x"0000";
    tmp(16072) := x"0000";
    tmp(16073) := x"0000";
    tmp(16074) := x"0000";
    tmp(16075) := x"0000";
    tmp(16076) := x"0000";
    tmp(16077) := x"0820";
    tmp(16078) := x"0820";
    tmp(16079) := x"0820";
    tmp(16080) := x"1040";
    tmp(16081) := x"bac0";
    tmp(16082) := x"b2a0";
    tmp(16083) := x"b2a0";
    tmp(16084) := x"baa0";
    tmp(16085) := x"baa0";
    tmp(16086) := x"baa0";
    tmp(16087) := x"bac0";
    tmp(16088) := x"c2c0";
    tmp(16089) := x"c2c0";
    tmp(16090) := x"cb00";
    tmp(16091) := x"cb20";
    tmp(16092) := x"c300";
    tmp(16093) := x"cb40";
    tmp(16094) := x"cb20";
    tmp(16095) := x"c2c0";
    tmp(16096) := x"c2e0";
    tmp(16097) := x"cb00";
    tmp(16098) := x"cb00";
    tmp(16099) := x"d320";
    tmp(16100) := x"db40";
    tmp(16101) := x"e340";
    tmp(16102) := x"db20";
    tmp(16103) := x"db00";
    tmp(16104) := x"db20";
    tmp(16105) := x"d320";
    tmp(16106) := x"db40";
    tmp(16107) := x"eb80";
    tmp(16108) := x"eba0";
    tmp(16109) := x"f3c0";
    tmp(16110) := x"eba0";
    tmp(16111) := x"fbe0";
    tmp(16112) := x"fc00";
    tmp(16113) := x"fc00";
    tmp(16114) := x"f440";
    tmp(16115) := x"f460";
    tmp(16116) := x"ec20";
    tmp(16117) := x"d360";
    tmp(16118) := x"bac0";
    tmp(16119) := x"a260";
    tmp(16120) := x"a240";
    tmp(16121) := x"a260";
    tmp(16122) := x"aaa0";
    tmp(16123) := x"aac0";
    tmp(16124) := x"b2c0";
    tmp(16125) := x"b2a0";
    tmp(16126) := x"b280";
    tmp(16127) := x"ba80";
    tmp(16128) := x"aa60";
    tmp(16129) := x"a220";
    tmp(16130) := x"9a00";
    tmp(16131) := x"9a00";
    tmp(16132) := x"91e0";
    tmp(16133) := x"89e0";
    tmp(16134) := x"89e0";
    tmp(16135) := x"9200";
    tmp(16136) := x"9a20";
    tmp(16137) := x"aa60";
    tmp(16138) := x"aa60";
    tmp(16139) := x"b260";
    tmp(16140) := x"b280";
    tmp(16141) := x"b280";
    tmp(16142) := x"aa40";
    tmp(16143) := x"9200";
    tmp(16144) := x"89c0";
    tmp(16145) := x"71a0";
    tmp(16146) := x"6160";
    tmp(16147) := x"4120";
    tmp(16148) := x"28c0";
    tmp(16149) := x"18a0";
    tmp(16150) := x"0840";
    tmp(16151) := x"0020";
    tmp(16152) := x"0000";
    tmp(16153) := x"0000";
    tmp(16154) := x"0020";
    tmp(16155) := x"0000";
    tmp(16156) := x"0000";
    tmp(16157) := x"0000";
    tmp(16158) := x"0000";
    tmp(16159) := x"0000";
    tmp(16160) := x"0000";
    tmp(16161) := x"0000";
    tmp(16162) := x"0000";
    tmp(16163) := x"0000";
    tmp(16164) := x"0000";
    tmp(16165) := x"0000";
    tmp(16166) := x"0000";
    tmp(16167) := x"0000";
    tmp(16168) := x"0000";
    tmp(16169) := x"0000";
    tmp(16170) := x"0000";
    tmp(16171) := x"0000";
    tmp(16172) := x"0000";
    tmp(16173) := x"0841";
    tmp(16174) := x"4185";
    tmp(16175) := x"6249";
    tmp(16176) := x"7acc";
    tmp(16177) := x"934f";
    tmp(16178) := x"a3f2";
    tmp(16179) := x"934f";
    tmp(16180) := x"c4b5";
    tmp(16181) := x"a3b0";
    tmp(16182) := x"bc52";
    tmp(16183) := x"934f";
    tmp(16184) := x"9b91";
    tmp(16185) := x"ac35";
    tmp(16186) := x"a3d2";
    tmp(16187) := x"9b4f";
    tmp(16188) := x"828c";
    tmp(16189) := x"ab90";
    tmp(16190) := x"c476";
    tmp(16191) := x"ccf7";
    tmp(16192) := x"fe9d";
    tmp(16193) := x"f5da";
    tmp(16194) := x"f5fb";
    tmp(16195) := x"ff3e";
    tmp(16196) := x"ed79";
    tmp(16197) := x"ff3d";
    tmp(16198) := x"ff1d";
    tmp(16199) := x"936d";
    tmp(16200) := x"0000";
    tmp(16201) := x"0000";
    tmp(16202) := x"49c6";
    tmp(16203) := x"ff1b";
    tmp(16204) := x"5a69";
    tmp(16205) := x"0820";
    tmp(16206) := x"49a6";
    tmp(16207) := x"c4f4";
    tmp(16208) := x"1082";
    tmp(16209) := x"18a2";
    tmp(16210) := x"72ab";
    tmp(16211) := x"93d0";
    tmp(16212) := x"0841";
    tmp(16213) := x"41a7";
    tmp(16214) := x"28e4";
    tmp(16215) := x"e61b";
    tmp(16216) := x"b4f5";
    tmp(16217) := x"7b2d";
    tmp(16218) := x"3985";
    tmp(16219) := x"0841";
    tmp(16220) := x"0841";
    tmp(16221) := x"1061";
    tmp(16222) := x"3165";
    tmp(16223) := x"31a5";
    tmp(16224) := x"0840";
    tmp(16225) := x"0880";
    tmp(16226) := x"08c0";
    tmp(16227) := x"10e0";
    tmp(16228) := x"10c0";
    tmp(16229) := x"1100";
    tmp(16230) := x"1940";
    tmp(16231) := x"1940";
    tmp(16232) := x"1960";
    tmp(16233) := x"21e0";
    tmp(16234) := x"19a0";
    tmp(16235) := x"21e0";
    tmp(16236) := x"3322";
    tmp(16237) := x"1161";
    tmp(16238) := x"0880";
    tmp(16239) := x"08a0";
    tmp(16240) := x"08a0";
    tmp(16241) := x"08a0";
    tmp(16242) := x"10c0";
    tmp(16243) := x"10c0";
    tmp(16244) := x"10e0";
    tmp(16245) := x"1100";
    tmp(16246) := x"1100";
    tmp(16247) := x"1100";
    tmp(16248) := x"1100";
    tmp(16249) := x"1100";
    tmp(16250) := x"1120";
    tmp(16251) := x"1120";
    tmp(16252) := x"1120";
    tmp(16253) := x"1120";
    tmp(16254) := x"1120";
    tmp(16255) := x"1100";
    tmp(16256) := x"0900";
    tmp(16257) := x"0900";
    tmp(16258) := x"08e0";
    tmp(16259) := x"08a0";
    tmp(16260) := x"08a0";
    tmp(16261) := x"08a0";
    tmp(16262) := x"0880";
    tmp(16263) := x"0880";
    tmp(16264) := x"0880";
    tmp(16265) := x"0860";
    tmp(16266) := x"0860";
    tmp(16267) := x"0860";
    tmp(16268) := x"0860";
    tmp(16269) := x"0860";
    tmp(16270) := x"0840";
    tmp(16271) := x"0840";
    tmp(16272) := x"0840";
    tmp(16273) := x"0840";
    tmp(16274) := x"0840";
    tmp(16275) := x"0820";
    tmp(16276) := x"0820";
    tmp(16277) := x"0000";
    tmp(16278) := x"0000";
    tmp(16279) := x"0000";
    tmp(16280) := x"0000";
    tmp(16281) := x"0000";
    tmp(16282) := x"0000";
    tmp(16283) := x"0000";
    tmp(16284) := x"0000";
    tmp(16285) := x"0000";
    tmp(16286) := x"0000";
    tmp(16287) := x"0000";
    tmp(16288) := x"0000";
    tmp(16289) := x"0000";
    tmp(16290) := x"0000";
    tmp(16291) := x"0000";
    tmp(16292) := x"0000";
    tmp(16293) := x"0000";
    tmp(16294) := x"0000";
    tmp(16295) := x"0000";
    tmp(16296) := x"0000";
    tmp(16297) := x"0000";
    tmp(16298) := x"0000";
    tmp(16299) := x"0000";
    tmp(16300) := x"0000";
    tmp(16301) := x"0000";
    tmp(16302) := x"0000";
    tmp(16303) := x"0000";
    tmp(16304) := x"0000";
    tmp(16305) := x"0000";
    tmp(16306) := x"0000";
    tmp(16307) := x"0000";
    tmp(16308) := x"0000";
    tmp(16309) := x"0000";
    tmp(16310) := x"0000";
    tmp(16311) := x"0000";
    tmp(16312) := x"0000";
    tmp(16313) := x"0000";
    tmp(16314) := x"0000";
    tmp(16315) := x"0000";
    tmp(16316) := x"0000";
    tmp(16317) := x"0820";
    tmp(16318) := x"0820";
    tmp(16319) := x"0820";
    tmp(16320) := x"1040";
    tmp(16321) := x"bac0";
    tmp(16322) := x"baa0";
    tmp(16323) := x"baa0";
    tmp(16324) := x"b2a0";
    tmp(16325) := x"b2c0";
    tmp(16326) := x"b2a0";
    tmp(16327) := x"bac0";
    tmp(16328) := x"c2e0";
    tmp(16329) := x"cb20";
    tmp(16330) := x"cb40";
    tmp(16331) := x"cb40";
    tmp(16332) := x"c320";
    tmp(16333) := x"d340";
    tmp(16334) := x"cb20";
    tmp(16335) := x"baa0";
    tmp(16336) := x"cac0";
    tmp(16337) := x"cae0";
    tmp(16338) := x"cae0";
    tmp(16339) := x"db20";
    tmp(16340) := x"cb00";
    tmp(16341) := x"d300";
    tmp(16342) := x"d2e0";
    tmp(16343) := x"d2e0";
    tmp(16344) := x"d300";
    tmp(16345) := x"d300";
    tmp(16346) := x"db20";
    tmp(16347) := x"db60";
    tmp(16348) := x"f3a0";
    tmp(16349) := x"fbe0";
    tmp(16350) := x"fc00";
    tmp(16351) := x"fc40";
    tmp(16352) := x"fc60";
    tmp(16353) := x"fcc0";
    tmp(16354) := x"fcc0";
    tmp(16355) := x"fcc0";
    tmp(16356) := x"f460";
    tmp(16357) := x"dba0";
    tmp(16358) := x"bae0";
    tmp(16359) := x"aa60";
    tmp(16360) := x"a240";
    tmp(16361) := x"a280";
    tmp(16362) := x"aaa0";
    tmp(16363) := x"aa80";
    tmp(16364) := x"aa80";
    tmp(16365) := x"b280";
    tmp(16366) := x"aa60";
    tmp(16367) := x"b260";
    tmp(16368) := x"b280";
    tmp(16369) := x"b280";
    tmp(16370) := x"aa60";
    tmp(16371) := x"9a00";
    tmp(16372) := x"91c0";
    tmp(16373) := x"91e0";
    tmp(16374) := x"9200";
    tmp(16375) := x"9200";
    tmp(16376) := x"a240";
    tmp(16377) := x"a220";
    tmp(16378) := x"aa40";
    tmp(16379) := x"b260";
    tmp(16380) := x"b260";
    tmp(16381) := x"b280";
    tmp(16382) := x"b260";
    tmp(16383) := x"91e0";
    tmp(16384) := x"81c0";
    tmp(16385) := x"7180";
    tmp(16386) := x"5940";
    tmp(16387) := x"4120";
    tmp(16388) := x"28c0";
    tmp(16389) := x"1080";
    tmp(16390) := x"0840";
    tmp(16391) := x"0020";
    tmp(16392) := x"0000";
    tmp(16393) := x"0020";
    tmp(16394) := x"0020";
    tmp(16395) := x"0000";
    tmp(16396) := x"0000";
    tmp(16397) := x"0000";
    tmp(16398) := x"0000";
    tmp(16399) := x"0000";
    tmp(16400) := x"0000";
    tmp(16401) := x"0000";
    tmp(16402) := x"0000";
    tmp(16403) := x"0000";
    tmp(16404) := x"0000";
    tmp(16405) := x"0000";
    tmp(16406) := x"0000";
    tmp(16407) := x"0000";
    tmp(16408) := x"0000";
    tmp(16409) := x"0000";
    tmp(16410) := x"0000";
    tmp(16411) := x"0000";
    tmp(16412) := x"0000";
    tmp(16413) := x"18a2";
    tmp(16414) := x"4185";
    tmp(16415) := x"6a4a";
    tmp(16416) := x"728b";
    tmp(16417) := x"8b2e";
    tmp(16418) := x"9bb1";
    tmp(16419) := x"934f";
    tmp(16420) := x"ddb9";
    tmp(16421) := x"c4b5";
    tmp(16422) := x"ddb8";
    tmp(16423) := x"c4d6";
    tmp(16424) := x"934f";
    tmp(16425) := x"b3f3";
    tmp(16426) := x"b413";
    tmp(16427) := x"bc33";
    tmp(16428) := x"7a4a";
    tmp(16429) := x"bbd2";
    tmp(16430) := x"b3d2";
    tmp(16431) := x"d4b5";
    tmp(16432) := x"ed37";
    tmp(16433) := x"ed98";
    tmp(16434) := x"fe9d";
    tmp(16435) := x"ed99";
    tmp(16436) := x"f69d";
    tmp(16437) := x"ffdf";
    tmp(16438) := x"ffdf";
    tmp(16439) := x"0841";
    tmp(16440) := x"0000";
    tmp(16441) := x"1041";
    tmp(16442) := x"feb9";
    tmp(16443) := x"cdf8";
    tmp(16444) := x"18a2";
    tmp(16445) := x"1861";
    tmp(16446) := x"ccd3";
    tmp(16447) := x"6a8a";
    tmp(16448) := x"1061";
    tmp(16449) := x"5228";
    tmp(16450) := x"3125";
    tmp(16451) := x"3966";
    tmp(16452) := x"2903";
    tmp(16453) := x"838d";
    tmp(16454) := x"0841";
    tmp(16455) := x"20a3";
    tmp(16456) := x"834f";
    tmp(16457) := x"b4f6";
    tmp(16458) := x"b4f4";
    tmp(16459) := x"a4b2";
    tmp(16460) := x"3185";
    tmp(16461) := x"0820";
    tmp(16462) := x"0820";
    tmp(16463) := x"18e2";
    tmp(16464) := x"0880";
    tmp(16465) := x"0880";
    tmp(16466) := x"08a0";
    tmp(16467) := x"08a0";
    tmp(16468) := x"08a0";
    tmp(16469) := x"1100";
    tmp(16470) := x"1920";
    tmp(16471) := x"1980";
    tmp(16472) := x"2180";
    tmp(16473) := x"21c0";
    tmp(16474) := x"19a0";
    tmp(16475) := x"2a81";
    tmp(16476) := x"3342";
    tmp(16477) := x"1120";
    tmp(16478) := x"0860";
    tmp(16479) := x"08a0";
    tmp(16480) := x"08a0";
    tmp(16481) := x"10c0";
    tmp(16482) := x"10c0";
    tmp(16483) := x"10e0";
    tmp(16484) := x"10e0";
    tmp(16485) := x"1100";
    tmp(16486) := x"1120";
    tmp(16487) := x"1120";
    tmp(16488) := x"1120";
    tmp(16489) := x"1120";
    tmp(16490) := x"1940";
    tmp(16491) := x"1940";
    tmp(16492) := x"1940";
    tmp(16493) := x"1960";
    tmp(16494) := x"1160";
    tmp(16495) := x"1140";
    tmp(16496) := x"1120";
    tmp(16497) := x"1120";
    tmp(16498) := x"0900";
    tmp(16499) := x"08e0";
    tmp(16500) := x"08c0";
    tmp(16501) := x"08c0";
    tmp(16502) := x"08a0";
    tmp(16503) := x"08a0";
    tmp(16504) := x"0880";
    tmp(16505) := x"0880";
    tmp(16506) := x"0860";
    tmp(16507) := x"0860";
    tmp(16508) := x"0860";
    tmp(16509) := x"0860";
    tmp(16510) := x"0840";
    tmp(16511) := x"0840";
    tmp(16512) := x"0840";
    tmp(16513) := x"0840";
    tmp(16514) := x"0840";
    tmp(16515) := x"0820";
    tmp(16516) := x"0820";
    tmp(16517) := x"0000";
    tmp(16518) := x"0000";
    tmp(16519) := x"0000";
    tmp(16520) := x"0000";
    tmp(16521) := x"0000";
    tmp(16522) := x"0000";
    tmp(16523) := x"0000";
    tmp(16524) := x"0000";
    tmp(16525) := x"0000";
    tmp(16526) := x"0000";
    tmp(16527) := x"0000";
    tmp(16528) := x"0000";
    tmp(16529) := x"0000";
    tmp(16530) := x"0000";
    tmp(16531) := x"0000";
    tmp(16532) := x"0000";
    tmp(16533) := x"0000";
    tmp(16534) := x"0000";
    tmp(16535) := x"0000";
    tmp(16536) := x"0000";
    tmp(16537) := x"0000";
    tmp(16538) := x"0000";
    tmp(16539) := x"0000";
    tmp(16540) := x"0000";
    tmp(16541) := x"0000";
    tmp(16542) := x"0000";
    tmp(16543) := x"0000";
    tmp(16544) := x"0000";
    tmp(16545) := x"0000";
    tmp(16546) := x"0000";
    tmp(16547) := x"0000";
    tmp(16548) := x"0000";
    tmp(16549) := x"0000";
    tmp(16550) := x"0000";
    tmp(16551) := x"0000";
    tmp(16552) := x"0000";
    tmp(16553) := x"0000";
    tmp(16554) := x"0000";
    tmp(16555) := x"0000";
    tmp(16556) := x"0000";
    tmp(16557) := x"0820";
    tmp(16558) := x"0820";
    tmp(16559) := x"0820";
    tmp(16560) := x"1040";
    tmp(16561) := x"bac0";
    tmp(16562) := x"b280";
    tmp(16563) := x"b280";
    tmp(16564) := x"b2a0";
    tmp(16565) := x"b2c0";
    tmp(16566) := x"bac0";
    tmp(16567) := x"bac0";
    tmp(16568) := x"bac0";
    tmp(16569) := x"cb20";
    tmp(16570) := x"cb40";
    tmp(16571) := x"cb40";
    tmp(16572) := x"d360";
    tmp(16573) := x"d360";
    tmp(16574) := x"d340";
    tmp(16575) := x"db60";
    tmp(16576) := x"d300";
    tmp(16577) := x"cac0";
    tmp(16578) := x"d320";
    tmp(16579) := x"db20";
    tmp(16580) := x"d300";
    tmp(16581) := x"db20";
    tmp(16582) := x"e340";
    tmp(16583) := x"cb00";
    tmp(16584) := x"cae0";
    tmp(16585) := x"cae0";
    tmp(16586) := x"db40";
    tmp(16587) := x"e380";
    tmp(16588) := x"eb80";
    tmp(16589) := x"f3c0";
    tmp(16590) := x"fc40";
    tmp(16591) := x"fc60";
    tmp(16592) := x"fc80";
    tmp(16593) := x"fd00";
    tmp(16594) := x"fd60";
    tmp(16595) := x"fd61";
    tmp(16596) := x"fd00";
    tmp(16597) := x"ec40";
    tmp(16598) := x"c320";
    tmp(16599) := x"aa80";
    tmp(16600) := x"a260";
    tmp(16601) := x"a260";
    tmp(16602) := x"aa80";
    tmp(16603) := x"aa80";
    tmp(16604) := x"aa80";
    tmp(16605) := x"a240";
    tmp(16606) := x"aa40";
    tmp(16607) := x"ba80";
    tmp(16608) := x"baa0";
    tmp(16609) := x"baa0";
    tmp(16610) := x"ba80";
    tmp(16611) := x"a220";
    tmp(16612) := x"9a00";
    tmp(16613) := x"9a20";
    tmp(16614) := x"9a00";
    tmp(16615) := x"a220";
    tmp(16616) := x"aa60";
    tmp(16617) := x"b260";
    tmp(16618) := x"ba80";
    tmp(16619) := x"b260";
    tmp(16620) := x"ba80";
    tmp(16621) := x"b260";
    tmp(16622) := x"aa40";
    tmp(16623) := x"9200";
    tmp(16624) := x"89e0";
    tmp(16625) := x"7180";
    tmp(16626) := x"5940";
    tmp(16627) := x"4100";
    tmp(16628) := x"20c0";
    tmp(16629) := x"1080";
    tmp(16630) := x"0860";
    tmp(16631) := x"0020";
    tmp(16632) := x"0000";
    tmp(16633) := x"0020";
    tmp(16634) := x"0020";
    tmp(16635) := x"0020";
    tmp(16636) := x"0000";
    tmp(16637) := x"0000";
    tmp(16638) := x"0000";
    tmp(16639) := x"0000";
    tmp(16640) := x"0000";
    tmp(16641) := x"0000";
    tmp(16642) := x"0000";
    tmp(16643) := x"0000";
    tmp(16644) := x"0000";
    tmp(16645) := x"0000";
    tmp(16646) := x"0000";
    tmp(16647) := x"0000";
    tmp(16648) := x"0000";
    tmp(16649) := x"0000";
    tmp(16650) := x"0000";
    tmp(16651) := x"0000";
    tmp(16652) := x"0000";
    tmp(16653) := x"2904";
    tmp(16654) := x"51c7";
    tmp(16655) := x"6229";
    tmp(16656) := x"728b";
    tmp(16657) := x"8b0e";
    tmp(16658) := x"936f";
    tmp(16659) := x"bc95";
    tmp(16660) := x"ccf7";
    tmp(16661) := x"edba";
    tmp(16662) := x"e5ba";
    tmp(16663) := x"fe3d";
    tmp(16664) := x"ccd6";
    tmp(16665) := x"b3b1";
    tmp(16666) := x"dcd7";
    tmp(16667) := x"8aee";
    tmp(16668) := x"ab6f";
    tmp(16669) := x"8acd";
    tmp(16670) := x"b3b2";
    tmp(16671) := x"b3b2";
    tmp(16672) := x"d454";
    tmp(16673) := x"f5b9";
    tmp(16674) := x"fe5c";
    tmp(16675) := x"ee3a";
    tmp(16676) := x"fe9b";
    tmp(16677) := x"ffff";
    tmp(16678) := x"41c7";
    tmp(16679) := x"0000";
    tmp(16680) := x"0000";
    tmp(16681) := x"938d";
    tmp(16682) := x"f69b";
    tmp(16683) := x"7b8e";
    tmp(16684) := x"0820";
    tmp(16685) := x"72ca";
    tmp(16686) := x"c4d3";
    tmp(16687) := x"20c3";
    tmp(16688) := x"1041";
    tmp(16689) := x"8b8e";
    tmp(16690) := x"20a3";
    tmp(16691) := x"2904";
    tmp(16692) := x"28e3";
    tmp(16693) := x"6aec";
    tmp(16694) := x"a472";
    tmp(16695) := x"0820";
    tmp(16696) := x"0821";
    tmp(16697) := x"20c4";
    tmp(16698) := x"2905";
    tmp(16699) := x"838f";
    tmp(16700) := x"18a3";
    tmp(16701) := x"83ad";
    tmp(16702) := x"39a5";
    tmp(16703) := x"0861";
    tmp(16704) := x"0860";
    tmp(16705) := x"0880";
    tmp(16706) := x"08a0";
    tmp(16707) := x"10e0";
    tmp(16708) := x"10e0";
    tmp(16709) := x"1120";
    tmp(16710) := x"1920";
    tmp(16711) := x"1940";
    tmp(16712) := x"1981";
    tmp(16713) := x"21a1";
    tmp(16714) := x"19c1";
    tmp(16715) := x"33a2";
    tmp(16716) := x"3342";
    tmp(16717) := x"08c0";
    tmp(16718) := x"0880";
    tmp(16719) := x"08a0";
    tmp(16720) := x"08a0";
    tmp(16721) := x"08c0";
    tmp(16722) := x"10c0";
    tmp(16723) := x"10e0";
    tmp(16724) := x"10e0";
    tmp(16725) := x"1900";
    tmp(16726) := x"1920";
    tmp(16727) := x"1940";
    tmp(16728) := x"1940";
    tmp(16729) := x"1940";
    tmp(16730) := x"1960";
    tmp(16731) := x"1961";
    tmp(16732) := x"1960";
    tmp(16733) := x"1960";
    tmp(16734) := x"1960";
    tmp(16735) := x"1960";
    tmp(16736) := x"1140";
    tmp(16737) := x"1140";
    tmp(16738) := x"1120";
    tmp(16739) := x"1120";
    tmp(16740) := x"1100";
    tmp(16741) := x"08e0";
    tmp(16742) := x"08c0";
    tmp(16743) := x"08a0";
    tmp(16744) := x"08a0";
    tmp(16745) := x"0880";
    tmp(16746) := x"0880";
    tmp(16747) := x"0880";
    tmp(16748) := x"0860";
    tmp(16749) := x"0860";
    tmp(16750) := x"0860";
    tmp(16751) := x"0860";
    tmp(16752) := x"0840";
    tmp(16753) := x"0840";
    tmp(16754) := x"0840";
    tmp(16755) := x"0840";
    tmp(16756) := x"0840";
    tmp(16757) := x"0000";
    tmp(16758) := x"0000";
    tmp(16759) := x"0000";
    tmp(16760) := x"0000";
    tmp(16761) := x"0000";
    tmp(16762) := x"0000";
    tmp(16763) := x"0000";
    tmp(16764) := x"0000";
    tmp(16765) := x"0000";
    tmp(16766) := x"0000";
    tmp(16767) := x"0000";
    tmp(16768) := x"0000";
    tmp(16769) := x"0000";
    tmp(16770) := x"0000";
    tmp(16771) := x"0000";
    tmp(16772) := x"0000";
    tmp(16773) := x"0000";
    tmp(16774) := x"0000";
    tmp(16775) := x"0000";
    tmp(16776) := x"0000";
    tmp(16777) := x"0000";
    tmp(16778) := x"0000";
    tmp(16779) := x"0000";
    tmp(16780) := x"0000";
    tmp(16781) := x"0000";
    tmp(16782) := x"0000";
    tmp(16783) := x"0000";
    tmp(16784) := x"0000";
    tmp(16785) := x"0000";
    tmp(16786) := x"0000";
    tmp(16787) := x"0000";
    tmp(16788) := x"0000";
    tmp(16789) := x"0000";
    tmp(16790) := x"0000";
    tmp(16791) := x"0000";
    tmp(16792) := x"0000";
    tmp(16793) := x"0000";
    tmp(16794) := x"0000";
    tmp(16795) := x"0000";
    tmp(16796) := x"0000";
    tmp(16797) := x"0820";
    tmp(16798) := x"0820";
    tmp(16799) := x"0820";
    tmp(16800) := x"1040";
    tmp(16801) := x"b280";
    tmp(16802) := x"aa60";
    tmp(16803) := x"b280";
    tmp(16804) := x"b2a0";
    tmp(16805) := x"bac0";
    tmp(16806) := x"b2c0";
    tmp(16807) := x"baa0";
    tmp(16808) := x"c2e0";
    tmp(16809) := x"cb40";
    tmp(16810) := x"cb40";
    tmp(16811) := x"cb00";
    tmp(16812) := x"cb20";
    tmp(16813) := x"d340";
    tmp(16814) := x"cb40";
    tmp(16815) := x"e360";
    tmp(16816) := x"d300";
    tmp(16817) := x"cb00";
    tmp(16818) := x"cae0";
    tmp(16819) := x"d300";
    tmp(16820) := x"d320";
    tmp(16821) := x"db20";
    tmp(16822) := x"db20";
    tmp(16823) := x"db40";
    tmp(16824) := x"db20";
    tmp(16825) := x"db40";
    tmp(16826) := x"db40";
    tmp(16827) := x"e340";
    tmp(16828) := x"eba0";
    tmp(16829) := x"f3c0";
    tmp(16830) := x"f3e0";
    tmp(16831) := x"fc00";
    tmp(16832) := x"fc60";
    tmp(16833) := x"fcc0";
    tmp(16834) := x"fd20";
    tmp(16835) := x"fd80";
    tmp(16836) := x"fd60";
    tmp(16837) := x"ec40";
    tmp(16838) := x"cb20";
    tmp(16839) := x"b2a0";
    tmp(16840) := x"aa60";
    tmp(16841) := x"aa80";
    tmp(16842) := x"aa80";
    tmp(16843) := x"aa60";
    tmp(16844) := x"aa60";
    tmp(16845) := x"aa60";
    tmp(16846) := x"b260";
    tmp(16847) := x"b260";
    tmp(16848) := x"b280";
    tmp(16849) := x"b2a0";
    tmp(16850) := x"b280";
    tmp(16851) := x"b260";
    tmp(16852) := x"9a00";
    tmp(16853) := x"91e0";
    tmp(16854) := x"9a20";
    tmp(16855) := x"a220";
    tmp(16856) := x"aa40";
    tmp(16857) := x"aa40";
    tmp(16858) := x"b260";
    tmp(16859) := x"b260";
    tmp(16860) := x"b260";
    tmp(16861) := x"b280";
    tmp(16862) := x"a240";
    tmp(16863) := x"9a20";
    tmp(16864) := x"9200";
    tmp(16865) := x"7180";
    tmp(16866) := x"5120";
    tmp(16867) := x"3900";
    tmp(16868) := x"20c0";
    tmp(16869) := x"1080";
    tmp(16870) := x"0840";
    tmp(16871) := x"0020";
    tmp(16872) := x"0000";
    tmp(16873) := x"0000";
    tmp(16874) := x"0020";
    tmp(16875) := x"0000";
    tmp(16876) := x"0000";
    tmp(16877) := x"0000";
    tmp(16878) := x"0000";
    tmp(16879) := x"0000";
    tmp(16880) := x"0000";
    tmp(16881) := x"0000";
    tmp(16882) := x"0000";
    tmp(16883) := x"0000";
    tmp(16884) := x"0000";
    tmp(16885) := x"0000";
    tmp(16886) := x"0000";
    tmp(16887) := x"0000";
    tmp(16888) := x"0000";
    tmp(16889) := x"0000";
    tmp(16890) := x"0000";
    tmp(16891) := x"0000";
    tmp(16892) := x"0820";
    tmp(16893) := x"41c7";
    tmp(16894) := x"49a7";
    tmp(16895) := x"6229";
    tmp(16896) := x"7acc";
    tmp(16897) := x"8b0e";
    tmp(16898) := x"9b90";
    tmp(16899) := x"abf2";
    tmp(16900) := x"d518";
    tmp(16901) := x"e579";
    tmp(16902) := x"f63b";
    tmp(16903) := x"fe7d";
    tmp(16904) := x"ff1f";
    tmp(16905) := x"c453";
    tmp(16906) := x"cc32";
    tmp(16907) := x"b3b0";
    tmp(16908) := x"930e";
    tmp(16909) := x"8aac";
    tmp(16910) := x"ab70";
    tmp(16911) := x"bbd1";
    tmp(16912) := x"dcf6";
    tmp(16913) := x"f5fb";
    tmp(16914) := x"fe3b";
    tmp(16915) := x"fe9c";
    tmp(16916) := x"ffdf";
    tmp(16917) := x"93f0";
    tmp(16918) := x"0000";
    tmp(16919) := x"0820";
    tmp(16920) := x"5a26";
    tmp(16921) := x"ccd3";
    tmp(16922) := x"bcd4";
    tmp(16923) := x"1041";
    tmp(16924) := x"28e3";
    tmp(16925) := x"d535";
    tmp(16926) := x"830c";
    tmp(16927) := x"0820";
    tmp(16928) := x"1081";
    tmp(16929) := x"9c31";
    tmp(16930) := x"28e4";
    tmp(16931) := x"5269";
    tmp(16932) := x"0841";
    tmp(16933) := x"5a6b";
    tmp(16934) := x"4188";
    tmp(16935) := x"8bcf";
    tmp(16936) := x"5a8a";
    tmp(16937) := x"0841";
    tmp(16938) := x"0821";
    tmp(16939) := x"2925";
    tmp(16940) := x"2945";
    tmp(16941) := x"1061";
    tmp(16942) := x"9c70";
    tmp(16943) := x"2102";
    tmp(16944) := x"0840";
    tmp(16945) := x"0880";
    tmp(16946) := x"08c0";
    tmp(16947) := x"08c0";
    tmp(16948) := x"1120";
    tmp(16949) := x"1120";
    tmp(16950) := x"1120";
    tmp(16951) := x"1960";
    tmp(16952) := x"1981";
    tmp(16953) := x"19c2";
    tmp(16954) := x"2262";
    tmp(16955) := x"3c03";
    tmp(16956) := x"2aa1";
    tmp(16957) := x"0880";
    tmp(16958) := x"0880";
    tmp(16959) := x"08a0";
    tmp(16960) := x"08a0";
    tmp(16961) := x"08a0";
    tmp(16962) := x"10c0";
    tmp(16963) := x"10e0";
    tmp(16964) := x"10e0";
    tmp(16965) := x"1921";
    tmp(16966) := x"1921";
    tmp(16967) := x"2161";
    tmp(16968) := x"2161";
    tmp(16969) := x"2161";
    tmp(16970) := x"2161";
    tmp(16971) := x"2161";
    tmp(16972) := x"2161";
    tmp(16973) := x"2161";
    tmp(16974) := x"1961";
    tmp(16975) := x"1960";
    tmp(16976) := x"1960";
    tmp(16977) := x"1960";
    tmp(16978) := x"1960";
    tmp(16979) := x"1160";
    tmp(16980) := x"1120";
    tmp(16981) := x"1120";
    tmp(16982) := x"1100";
    tmp(16983) := x"08e0";
    tmp(16984) := x"08c0";
    tmp(16985) := x"08a0";
    tmp(16986) := x"0880";
    tmp(16987) := x"0880";
    tmp(16988) := x"0880";
    tmp(16989) := x"0860";
    tmp(16990) := x"0860";
    tmp(16991) := x"0860";
    tmp(16992) := x"0860";
    tmp(16993) := x"0840";
    tmp(16994) := x"0840";
    tmp(16995) := x"0840";
    tmp(16996) := x"0840";
    tmp(16997) := x"0000";
    tmp(16998) := x"0000";
    tmp(16999) := x"0000";
    tmp(17000) := x"0000";
    tmp(17001) := x"0000";
    tmp(17002) := x"0000";
    tmp(17003) := x"0000";
    tmp(17004) := x"0000";
    tmp(17005) := x"0000";
    tmp(17006) := x"0000";
    tmp(17007) := x"0000";
    tmp(17008) := x"0000";
    tmp(17009) := x"0000";
    tmp(17010) := x"0000";
    tmp(17011) := x"0000";
    tmp(17012) := x"0000";
    tmp(17013) := x"0000";
    tmp(17014) := x"0000";
    tmp(17015) := x"0000";
    tmp(17016) := x"0000";
    tmp(17017) := x"0000";
    tmp(17018) := x"0000";
    tmp(17019) := x"0000";
    tmp(17020) := x"0000";
    tmp(17021) := x"0000";
    tmp(17022) := x"0000";
    tmp(17023) := x"0000";
    tmp(17024) := x"0000";
    tmp(17025) := x"0000";
    tmp(17026) := x"0000";
    tmp(17027) := x"0000";
    tmp(17028) := x"0000";
    tmp(17029) := x"0000";
    tmp(17030) := x"0000";
    tmp(17031) := x"0000";
    tmp(17032) := x"0000";
    tmp(17033) := x"0000";
    tmp(17034) := x"0000";
    tmp(17035) := x"0000";
    tmp(17036) := x"0000";
    tmp(17037) := x"0820";
    tmp(17038) := x"0820";
    tmp(17039) := x"0820";
    tmp(17040) := x"1040";
    tmp(17041) := x"aa80";
    tmp(17042) := x"a260";
    tmp(17043) := x"aa80";
    tmp(17044) := x"aa80";
    tmp(17045) := x"aa80";
    tmp(17046) := x"aa80";
    tmp(17047) := x"aa80";
    tmp(17048) := x"bac0";
    tmp(17049) := x"c2e0";
    tmp(17050) := x"c300";
    tmp(17051) := x"c320";
    tmp(17052) := x"cb20";
    tmp(17053) := x"cb40";
    tmp(17054) := x"d360";
    tmp(17055) := x"db60";
    tmp(17056) := x"eb60";
    tmp(17057) := x"d300";
    tmp(17058) := x"cb00";
    tmp(17059) := x"d2e0";
    tmp(17060) := x"d2e0";
    tmp(17061) := x"db20";
    tmp(17062) := x"e320";
    tmp(17063) := x"db20";
    tmp(17064) := x"db20";
    tmp(17065) := x"db40";
    tmp(17066) := x"db40";
    tmp(17067) := x"eb60";
    tmp(17068) := x"eb80";
    tmp(17069) := x"f3c0";
    tmp(17070) := x"fc00";
    tmp(17071) := x"fc00";
    tmp(17072) := x"fc40";
    tmp(17073) := x"fcc0";
    tmp(17074) := x"fd20";
    tmp(17075) := x"fd40";
    tmp(17076) := x"fca0";
    tmp(17077) := x"e380";
    tmp(17078) := x"c2c0";
    tmp(17079) := x"aa60";
    tmp(17080) := x"9a20";
    tmp(17081) := x"a260";
    tmp(17082) := x"aa60";
    tmp(17083) := x"aa60";
    tmp(17084) := x"ba80";
    tmp(17085) := x"b280";
    tmp(17086) := x"b280";
    tmp(17087) := x"b280";
    tmp(17088) := x"b280";
    tmp(17089) := x"bac0";
    tmp(17090) := x"baa0";
    tmp(17091) := x"b280";
    tmp(17092) := x"a240";
    tmp(17093) := x"9a20";
    tmp(17094) := x"9a00";
    tmp(17095) := x"9a20";
    tmp(17096) := x"aa40";
    tmp(17097) := x"b260";
    tmp(17098) := x"b260";
    tmp(17099) := x"b240";
    tmp(17100) := x"b260";
    tmp(17101) := x"aa60";
    tmp(17102) := x"aa60";
    tmp(17103) := x"a220";
    tmp(17104) := x"91e0";
    tmp(17105) := x"6980";
    tmp(17106) := x"5120";
    tmp(17107) := x"3900";
    tmp(17108) := x"20a0";
    tmp(17109) := x"1080";
    tmp(17110) := x"0860";
    tmp(17111) := x"0020";
    tmp(17112) := x"0020";
    tmp(17113) := x"0020";
    tmp(17114) := x"0000";
    tmp(17115) := x"0000";
    tmp(17116) := x"0000";
    tmp(17117) := x"0000";
    tmp(17118) := x"0000";
    tmp(17119) := x"0000";
    tmp(17120) := x"0000";
    tmp(17121) := x"0000";
    tmp(17122) := x"0000";
    tmp(17123) := x"0000";
    tmp(17124) := x"0000";
    tmp(17125) := x"0000";
    tmp(17126) := x"0000";
    tmp(17127) := x"0000";
    tmp(17128) := x"0000";
    tmp(17129) := x"0000";
    tmp(17130) := x"0000";
    tmp(17131) := x"0000";
    tmp(17132) := x"1061";
    tmp(17133) := x"3966";
    tmp(17134) := x"49c7";
    tmp(17135) := x"6228";
    tmp(17136) := x"7acc";
    tmp(17137) := x"8b0e";
    tmp(17138) := x"abd2";
    tmp(17139) := x"b413";
    tmp(17140) := x"dcf7";
    tmp(17141) := x"ed79";
    tmp(17142) := x"fe7d";
    tmp(17143) := x"f69c";
    tmp(17144) := x"ff9f";
    tmp(17145) := x"fe3c";
    tmp(17146) := x"d495";
    tmp(17147) := x"dc75";
    tmp(17148) := x"92cd";
    tmp(17149) := x"8a8c";
    tmp(17150) := x"92cc";
    tmp(17151) := x"bbb1";
    tmp(17152) := x"ed79";
    tmp(17153) := x"eddb";
    tmp(17154) := x"edb9";
    tmp(17155) := x"fe9b";
    tmp(17156) := x"ff9f";
    tmp(17157) := x"1061";
    tmp(17158) := x"0820";
    tmp(17159) := x"0841";
    tmp(17160) := x"ac0f";
    tmp(17161) := x"dd96";
    tmp(17162) := x"5a8a";
    tmp(17163) := x"0000";
    tmp(17164) := x"6a69";
    tmp(17165) := x"bc94";
    tmp(17166) := x"6aab";
    tmp(17167) := x"1061";
    tmp(17168) := x"3986";
    tmp(17169) := x"bcf6";
    tmp(17170) := x"41a7";
    tmp(17171) := x"4a08";
    tmp(17172) := x"3145";
    tmp(17173) := x"734e";
    tmp(17174) := x"49e8";
    tmp(17175) := x"2905";
    tmp(17176) := x"628b";
    tmp(17177) := x"cdf8";
    tmp(17178) := x"3185";
    tmp(17179) := x"0821";
    tmp(17180) := x"39a6";
    tmp(17181) := x"0841";
    tmp(17182) := x"3144";
    tmp(17183) := x"2142";
    tmp(17184) := x"0860";
    tmp(17185) := x"0880";
    tmp(17186) := x"08c0";
    tmp(17187) := x"10e0";
    tmp(17188) := x"1100";
    tmp(17189) := x"1100";
    tmp(17190) := x"1940";
    tmp(17191) := x"1940";
    tmp(17192) := x"1981";
    tmp(17193) := x"1981";
    tmp(17194) := x"2aa2";
    tmp(17195) := x"3ba1";
    tmp(17196) := x"19c0";
    tmp(17197) := x"0860";
    tmp(17198) := x"0880";
    tmp(17199) := x"08a0";
    tmp(17200) := x"08a0";
    tmp(17201) := x"08a0";
    tmp(17202) := x"10a0";
    tmp(17203) := x"10c0";
    tmp(17204) := x"1901";
    tmp(17205) := x"1921";
    tmp(17206) := x"2141";
    tmp(17207) := x"2141";
    tmp(17208) := x"2161";
    tmp(17209) := x"2981";
    tmp(17210) := x"2981";
    tmp(17211) := x"2161";
    tmp(17212) := x"2161";
    tmp(17213) := x"2161";
    tmp(17214) := x"2181";
    tmp(17215) := x"2181";
    tmp(17216) := x"1961";
    tmp(17217) := x"1981";
    tmp(17218) := x"1960";
    tmp(17219) := x"1960";
    tmp(17220) := x"1960";
    tmp(17221) := x"1940";
    tmp(17222) := x"1120";
    tmp(17223) := x"1100";
    tmp(17224) := x"1100";
    tmp(17225) := x"08e0";
    tmp(17226) := x"08c0";
    tmp(17227) := x"08a0";
    tmp(17228) := x"0880";
    tmp(17229) := x"0880";
    tmp(17230) := x"0860";
    tmp(17231) := x"0860";
    tmp(17232) := x"0860";
    tmp(17233) := x"0840";
    tmp(17234) := x"0840";
    tmp(17235) := x"0840";
    tmp(17236) := x"0840";
    tmp(17237) := x"0000";
    tmp(17238) := x"0000";
    tmp(17239) := x"0000";
    tmp(17240) := x"0000";
    tmp(17241) := x"0000";
    tmp(17242) := x"0000";
    tmp(17243) := x"0000";
    tmp(17244) := x"0000";
    tmp(17245) := x"0000";
    tmp(17246) := x"0000";
    tmp(17247) := x"0000";
    tmp(17248) := x"0000";
    tmp(17249) := x"0000";
    tmp(17250) := x"0000";
    tmp(17251) := x"0000";
    tmp(17252) := x"0000";
    tmp(17253) := x"0000";
    tmp(17254) := x"0000";
    tmp(17255) := x"0000";
    tmp(17256) := x"0000";
    tmp(17257) := x"0000";
    tmp(17258) := x"0000";
    tmp(17259) := x"0000";
    tmp(17260) := x"0000";
    tmp(17261) := x"0000";
    tmp(17262) := x"0000";
    tmp(17263) := x"0000";
    tmp(17264) := x"0000";
    tmp(17265) := x"0000";
    tmp(17266) := x"0000";
    tmp(17267) := x"0000";
    tmp(17268) := x"0000";
    tmp(17269) := x"0000";
    tmp(17270) := x"0000";
    tmp(17271) := x"0000";
    tmp(17272) := x"0000";
    tmp(17273) := x"0000";
    tmp(17274) := x"0000";
    tmp(17275) := x"0000";
    tmp(17276) := x"0000";
    tmp(17277) := x"0820";
    tmp(17278) := x"0820";
    tmp(17279) := x"0820";
    tmp(17280) := x"1040";
    tmp(17281) := x"b280";
    tmp(17282) := x"9a40";
    tmp(17283) := x"aa80";
    tmp(17284) := x"aa80";
    tmp(17285) := x"b280";
    tmp(17286) := x"aa60";
    tmp(17287) := x"aa60";
    tmp(17288) := x"b280";
    tmp(17289) := x"c2c0";
    tmp(17290) := x"d340";
    tmp(17291) := x"bac0";
    tmp(17292) := x"c300";
    tmp(17293) := x"cb20";
    tmp(17294) := x"d340";
    tmp(17295) := x"db40";
    tmp(17296) := x"d300";
    tmp(17297) := x"db20";
    tmp(17298) := x"db20";
    tmp(17299) := x"d2e0";
    tmp(17300) := x"dae0";
    tmp(17301) := x"db00";
    tmp(17302) := x"db00";
    tmp(17303) := x"d300";
    tmp(17304) := x"db20";
    tmp(17305) := x"e340";
    tmp(17306) := x"e340";
    tmp(17307) := x"eb60";
    tmp(17308) := x"eb60";
    tmp(17309) := x"fbe0";
    tmp(17310) := x"fc00";
    tmp(17311) := x"fc20";
    tmp(17312) := x"fc60";
    tmp(17313) := x"fca0";
    tmp(17314) := x"fd00";
    tmp(17315) := x"fce0";
    tmp(17316) := x"f400";
    tmp(17317) := x"db60";
    tmp(17318) := x"c2e0";
    tmp(17319) := x"c2a0";
    tmp(17320) := x"b260";
    tmp(17321) := x"aa60";
    tmp(17322) := x"b260";
    tmp(17323) := x"aa60";
    tmp(17324) := x"b280";
    tmp(17325) := x"b260";
    tmp(17326) := x"ba80";
    tmp(17327) := x"c280";
    tmp(17328) := x"baa0";
    tmp(17329) := x"baa0";
    tmp(17330) := x"baa0";
    tmp(17331) := x"aa40";
    tmp(17332) := x"a240";
    tmp(17333) := x"a220";
    tmp(17334) := x"aa40";
    tmp(17335) := x"aa60";
    tmp(17336) := x"b260";
    tmp(17337) := x"b260";
    tmp(17338) := x"b240";
    tmp(17339) := x"b240";
    tmp(17340) := x"aa40";
    tmp(17341) := x"aa40";
    tmp(17342) := x"aa40";
    tmp(17343) := x"a240";
    tmp(17344) := x"91e0";
    tmp(17345) := x"7180";
    tmp(17346) := x"5120";
    tmp(17347) := x"30e0";
    tmp(17348) := x"20a0";
    tmp(17349) := x"1080";
    tmp(17350) := x"0860";
    tmp(17351) := x"0020";
    tmp(17352) := x"0020";
    tmp(17353) := x"0000";
    tmp(17354) := x"0000";
    tmp(17355) := x"0000";
    tmp(17356) := x"0000";
    tmp(17357) := x"0000";
    tmp(17358) := x"0000";
    tmp(17359) := x"0000";
    tmp(17360) := x"0000";
    tmp(17361) := x"0000";
    tmp(17362) := x"0000";
    tmp(17363) := x"0000";
    tmp(17364) := x"0000";
    tmp(17365) := x"0000";
    tmp(17366) := x"0000";
    tmp(17367) := x"0000";
    tmp(17368) := x"0000";
    tmp(17369) := x"0000";
    tmp(17370) := x"0000";
    tmp(17371) := x"0000";
    tmp(17372) := x"0861";
    tmp(17373) := x"3986";
    tmp(17374) := x"51e8";
    tmp(17375) := x"59e8";
    tmp(17376) := x"7a6b";
    tmp(17377) := x"828c";
    tmp(17378) := x"a3b1";
    tmp(17379) := x"bc54";
    tmp(17380) := x"bc53";
    tmp(17381) := x"ed99";
    tmp(17382) := x"fede";
    tmp(17383) := x"ed78";
    tmp(17384) := x"ff1e";
    tmp(17385) := x"ff1f";
    tmp(17386) := x"f559";
    tmp(17387) := x"f5da";
    tmp(17388) := x"ab50";
    tmp(17389) := x"826b";
    tmp(17390) := x"928b";
    tmp(17391) := x"bbd0";
    tmp(17392) := x"ed38";
    tmp(17393) := x"ed79";
    tmp(17394) := x"ed99";
    tmp(17395) := x"ff9e";
    tmp(17396) := x"de39";
    tmp(17397) := x"2924";
    tmp(17398) := x"0000";
    tmp(17399) := x"0820";
    tmp(17400) := x"b471";
    tmp(17401) := x"e65a";
    tmp(17402) := x"1081";
    tmp(17403) := x"0841";
    tmp(17404) := x"e5d7";
    tmp(17405) := x"93b0";
    tmp(17406) := x"18a2";
    tmp(17407) := x"1061";
    tmp(17408) := x"7b4d";
    tmp(17409) := x"ac54";
    tmp(17410) := x"6aac";
    tmp(17411) := x"20a3";
    tmp(17412) := x"41c7";
    tmp(17413) := x"5a6b";
    tmp(17414) := x"acb4";
    tmp(17415) := x"2904";
    tmp(17416) := x"0841";
    tmp(17417) := x"3125";
    tmp(17418) := x"8bd0";
    tmp(17419) := x"2104";
    tmp(17420) := x"1061";
    tmp(17421) := x"41c6";
    tmp(17422) := x"18c2";
    tmp(17423) := x"0860";
    tmp(17424) := x"0860";
    tmp(17425) := x"08a0";
    tmp(17426) := x"08a0";
    tmp(17427) := x"10c0";
    tmp(17428) := x"10e0";
    tmp(17429) := x"1920";
    tmp(17430) := x"1120";
    tmp(17431) := x"1120";
    tmp(17432) := x"1981";
    tmp(17433) := x"19c1";
    tmp(17434) := x"2aa1";
    tmp(17435) := x"3321";
    tmp(17436) := x"08e0";
    tmp(17437) := x"0880";
    tmp(17438) := x"0880";
    tmp(17439) := x"08a0";
    tmp(17440) := x"08a0";
    tmp(17441) := x"08a0";
    tmp(17442) := x"10c0";
    tmp(17443) := x"10e0";
    tmp(17444) := x"1901";
    tmp(17445) := x"1921";
    tmp(17446) := x"2141";
    tmp(17447) := x"2141";
    tmp(17448) := x"2141";
    tmp(17449) := x"2981";
    tmp(17450) := x"2981";
    tmp(17451) := x"2981";
    tmp(17452) := x"2981";
    tmp(17453) := x"2981";
    tmp(17454) := x"2181";
    tmp(17455) := x"2161";
    tmp(17456) := x"2181";
    tmp(17457) := x"2181";
    tmp(17458) := x"2181";
    tmp(17459) := x"2161";
    tmp(17460) := x"1961";
    tmp(17461) := x"1960";
    tmp(17462) := x"1960";
    tmp(17463) := x"1120";
    tmp(17464) := x"1120";
    tmp(17465) := x"1100";
    tmp(17466) := x"08e0";
    tmp(17467) := x"08c0";
    tmp(17468) := x"08a0";
    tmp(17469) := x"08a0";
    tmp(17470) := x"0880";
    tmp(17471) := x"0860";
    tmp(17472) := x"0860";
    tmp(17473) := x"0860";
    tmp(17474) := x"0860";
    tmp(17475) := x"0840";
    tmp(17476) := x"0840";
    tmp(17477) := x"0000";
    tmp(17478) := x"0000";
    tmp(17479) := x"0000";
    tmp(17480) := x"0000";
    tmp(17481) := x"0000";
    tmp(17482) := x"0000";
    tmp(17483) := x"0000";
    tmp(17484) := x"0000";
    tmp(17485) := x"0000";
    tmp(17486) := x"0000";
    tmp(17487) := x"0000";
    tmp(17488) := x"0000";
    tmp(17489) := x"0000";
    tmp(17490) := x"0000";
    tmp(17491) := x"0000";
    tmp(17492) := x"0000";
    tmp(17493) := x"0000";
    tmp(17494) := x"0000";
    tmp(17495) := x"0000";
    tmp(17496) := x"0000";
    tmp(17497) := x"0000";
    tmp(17498) := x"0000";
    tmp(17499) := x"0000";
    tmp(17500) := x"0000";
    tmp(17501) := x"0000";
    tmp(17502) := x"0000";
    tmp(17503) := x"0000";
    tmp(17504) := x"0000";
    tmp(17505) := x"0000";
    tmp(17506) := x"0000";
    tmp(17507) := x"0000";
    tmp(17508) := x"0000";
    tmp(17509) := x"0000";
    tmp(17510) := x"0000";
    tmp(17511) := x"0000";
    tmp(17512) := x"0000";
    tmp(17513) := x"0000";
    tmp(17514) := x"0000";
    tmp(17515) := x"0000";
    tmp(17516) := x"0000";
    tmp(17517) := x"0820";
    tmp(17518) := x"0820";
    tmp(17519) := x"0840";
    tmp(17520) := x"1040";
    tmp(17521) := x"aa60";
    tmp(17522) := x"a260";
    tmp(17523) := x"a260";
    tmp(17524) := x"aa80";
    tmp(17525) := x"a280";
    tmp(17526) := x"aaa0";
    tmp(17527) := x"aa80";
    tmp(17528) := x"b280";
    tmp(17529) := x"b280";
    tmp(17530) := x"b2a0";
    tmp(17531) := x"bac0";
    tmp(17532) := x"c2e0";
    tmp(17533) := x"c2e0";
    tmp(17534) := x"cb40";
    tmp(17535) := x"d320";
    tmp(17536) := x"db20";
    tmp(17537) := x"db20";
    tmp(17538) := x"db00";
    tmp(17539) := x"cac0";
    tmp(17540) := x"d2e0";
    tmp(17541) := x"db00";
    tmp(17542) := x"e320";
    tmp(17543) := x"db40";
    tmp(17544) := x"e340";
    tmp(17545) := x"eb40";
    tmp(17546) := x"f360";
    tmp(17547) := x"eb40";
    tmp(17548) := x"f360";
    tmp(17549) := x"fbc0";
    tmp(17550) := x"fc00";
    tmp(17551) := x"fc00";
    tmp(17552) := x"fc40";
    tmp(17553) := x"fca0";
    tmp(17554) := x"fc80";
    tmp(17555) := x"fc40";
    tmp(17556) := x"f3c0";
    tmp(17557) := x"db60";
    tmp(17558) := x"cae0";
    tmp(17559) := x"c2a0";
    tmp(17560) := x"b280";
    tmp(17561) := x"b260";
    tmp(17562) := x"aa80";
    tmp(17563) := x"aa60";
    tmp(17564) := x"b280";
    tmp(17565) := x"b260";
    tmp(17566) := x"ba80";
    tmp(17567) := x"c280";
    tmp(17568) := x"b260";
    tmp(17569) := x"b280";
    tmp(17570) := x"b260";
    tmp(17571) := x"a240";
    tmp(17572) := x"9a20";
    tmp(17573) := x"9a20";
    tmp(17574) := x"a220";
    tmp(17575) := x"aa40";
    tmp(17576) := x"b260";
    tmp(17577) := x"b240";
    tmp(17578) := x"b240";
    tmp(17579) := x"b240";
    tmp(17580) := x"aa20";
    tmp(17581) := x"b240";
    tmp(17582) := x"aa40";
    tmp(17583) := x"a240";
    tmp(17584) := x"91e0";
    tmp(17585) := x"79a0";
    tmp(17586) := x"5940";
    tmp(17587) := x"4900";
    tmp(17588) := x"28c0";
    tmp(17589) := x"18a0";
    tmp(17590) := x"1080";
    tmp(17591) := x"0860";
    tmp(17592) := x"0020";
    tmp(17593) := x"0000";
    tmp(17594) := x"0000";
    tmp(17595) := x"0000";
    tmp(17596) := x"0000";
    tmp(17597) := x"0000";
    tmp(17598) := x"0000";
    tmp(17599) := x"0000";
    tmp(17600) := x"0000";
    tmp(17601) := x"0000";
    tmp(17602) := x"0000";
    tmp(17603) := x"0000";
    tmp(17604) := x"0000";
    tmp(17605) := x"0000";
    tmp(17606) := x"0000";
    tmp(17607) := x"0000";
    tmp(17608) := x"0000";
    tmp(17609) := x"0000";
    tmp(17610) := x"0000";
    tmp(17611) := x"0000";
    tmp(17612) := x"0821";
    tmp(17613) := x"2905";
    tmp(17614) := x"5209";
    tmp(17615) := x"59e8";
    tmp(17616) := x"6a09";
    tmp(17617) := x"92cd";
    tmp(17618) := x"930d";
    tmp(17619) := x"d495";
    tmp(17620) := x"bbf2";
    tmp(17621) := x"dcf6";
    tmp(17622) := x"f61a";
    tmp(17623) := x"ed99";
    tmp(17624) := x"fefd";
    tmp(17625) := x"ff1f";
    tmp(17626) := x"fdb9";
    tmp(17627) := x"ff1e";
    tmp(17628) := x"c3f3";
    tmp(17629) := x"8a8b";
    tmp(17630) := x"928b";
    tmp(17631) := x"bbaf";
    tmp(17632) := x"e4b5";
    tmp(17633) := x"ed38";
    tmp(17634) := x"e5b8";
    tmp(17635) := x"fedd";
    tmp(17636) := x"a492";
    tmp(17637) := x"0020";
    tmp(17638) := x"0000";
    tmp(17639) := x"1881";
    tmp(17640) := x"ee38";
    tmp(17641) := x"a451";
    tmp(17642) := x"0000";
    tmp(17643) := x"3985";
    tmp(17644) := x"e5b8";
    tmp(17645) := x"3125";
    tmp(17646) := x"0020";
    tmp(17647) := x"3965";
    tmp(17648) := x"a413";
    tmp(17649) := x"8b51";
    tmp(17650) := x"834f";
    tmp(17651) := x"524a";
    tmp(17652) := x"0821";
    tmp(17653) := x"6acc";
    tmp(17654) := x"18a3";
    tmp(17655) := x"6acc";
    tmp(17656) := x"732c";
    tmp(17657) := x"0000";
    tmp(17658) := x"0821";
    tmp(17659) := x"18c3";
    tmp(17660) := x"2924";
    tmp(17661) := x"3144";
    tmp(17662) := x"10a1";
    tmp(17663) := x"0040";
    tmp(17664) := x"0880";
    tmp(17665) := x"08c0";
    tmp(17666) := x"10c0";
    tmp(17667) := x"10c0";
    tmp(17668) := x"10e0";
    tmp(17669) := x"1100";
    tmp(17670) := x"10e0";
    tmp(17671) := x"1120";
    tmp(17672) := x"1980";
    tmp(17673) := x"2241";
    tmp(17674) := x"2ac1";
    tmp(17675) := x"2240";
    tmp(17676) := x"0880";
    tmp(17677) := x"0880";
    tmp(17678) := x"0880";
    tmp(17679) := x"08a0";
    tmp(17680) := x"08a0";
    tmp(17681) := x"08c0";
    tmp(17682) := x"10c0";
    tmp(17683) := x"10e0";
    tmp(17684) := x"1901";
    tmp(17685) := x"1901";
    tmp(17686) := x"2121";
    tmp(17687) := x"2141";
    tmp(17688) := x"2941";
    tmp(17689) := x"2961";
    tmp(17690) := x"2962";
    tmp(17691) := x"3182";
    tmp(17692) := x"31a2";
    tmp(17693) := x"2981";
    tmp(17694) := x"2981";
    tmp(17695) := x"2981";
    tmp(17696) := x"2161";
    tmp(17697) := x"2181";
    tmp(17698) := x"2181";
    tmp(17699) := x"2161";
    tmp(17700) := x"2161";
    tmp(17701) := x"2181";
    tmp(17702) := x"1961";
    tmp(17703) := x"1940";
    tmp(17704) := x"1940";
    tmp(17705) := x"1140";
    tmp(17706) := x"1100";
    tmp(17707) := x"1100";
    tmp(17708) := x"08e0";
    tmp(17709) := x"08a0";
    tmp(17710) := x"08a0";
    tmp(17711) := x"0880";
    tmp(17712) := x"0860";
    tmp(17713) := x"0860";
    tmp(17714) := x"0860";
    tmp(17715) := x"0860";
    tmp(17716) := x"0840";
    tmp(17717) := x"0000";
    tmp(17718) := x"0000";
    tmp(17719) := x"0000";
    tmp(17720) := x"0000";
    tmp(17721) := x"0000";
    tmp(17722) := x"0000";
    tmp(17723) := x"0000";
    tmp(17724) := x"0000";
    tmp(17725) := x"0000";
    tmp(17726) := x"0000";
    tmp(17727) := x"0000";
    tmp(17728) := x"0000";
    tmp(17729) := x"0000";
    tmp(17730) := x"0000";
    tmp(17731) := x"0000";
    tmp(17732) := x"0000";
    tmp(17733) := x"0000";
    tmp(17734) := x"0000";
    tmp(17735) := x"0000";
    tmp(17736) := x"0000";
    tmp(17737) := x"0000";
    tmp(17738) := x"0000";
    tmp(17739) := x"0000";
    tmp(17740) := x"0000";
    tmp(17741) := x"0000";
    tmp(17742) := x"0000";
    tmp(17743) := x"0000";
    tmp(17744) := x"0000";
    tmp(17745) := x"0000";
    tmp(17746) := x"0000";
    tmp(17747) := x"0000";
    tmp(17748) := x"0000";
    tmp(17749) := x"0000";
    tmp(17750) := x"0000";
    tmp(17751) := x"0000";
    tmp(17752) := x"0000";
    tmp(17753) := x"0000";
    tmp(17754) := x"0000";
    tmp(17755) := x"0000";
    tmp(17756) := x"0000";
    tmp(17757) := x"0820";
    tmp(17758) := x"0840";
    tmp(17759) := x"0840";
    tmp(17760) := x"1040";
    tmp(17761) := x"a240";
    tmp(17762) := x"9a40";
    tmp(17763) := x"a240";
    tmp(17764) := x"a260";
    tmp(17765) := x"aa60";
    tmp(17766) := x"aa80";
    tmp(17767) := x"b2a0";
    tmp(17768) := x"b280";
    tmp(17769) := x"b280";
    tmp(17770) := x"b2a0";
    tmp(17771) := x"bac0";
    tmp(17772) := x"c2e0";
    tmp(17773) := x"c2e0";
    tmp(17774) := x"cb20";
    tmp(17775) := x"d300";
    tmp(17776) := x"db40";
    tmp(17777) := x"db20";
    tmp(17778) := x"db00";
    tmp(17779) := x"d300";
    tmp(17780) := x"d300";
    tmp(17781) := x"e320";
    tmp(17782) := x"e320";
    tmp(17783) := x"eb40";
    tmp(17784) := x"eb60";
    tmp(17785) := x"eb60";
    tmp(17786) := x"f360";
    tmp(17787) := x"eb40";
    tmp(17788) := x"f380";
    tmp(17789) := x"fba0";
    tmp(17790) := x"fbe0";
    tmp(17791) := x"fc40";
    tmp(17792) := x"fc60";
    tmp(17793) := x"fc60";
    tmp(17794) := x"fc60";
    tmp(17795) := x"fc40";
    tmp(17796) := x"f3c0";
    tmp(17797) := x"e340";
    tmp(17798) := x"d300";
    tmp(17799) := x"c2a0";
    tmp(17800) := x"b260";
    tmp(17801) := x"aa60";
    tmp(17802) := x"aa40";
    tmp(17803) := x"aa20";
    tmp(17804) := x"b260";
    tmp(17805) := x"b260";
    tmp(17806) := x"b260";
    tmp(17807) := x"b280";
    tmp(17808) := x"b280";
    tmp(17809) := x"b280";
    tmp(17810) := x"a240";
    tmp(17811) := x"9a20";
    tmp(17812) := x"a220";
    tmp(17813) := x"aa20";
    tmp(17814) := x"aa40";
    tmp(17815) := x"aa40";
    tmp(17816) := x"ba80";
    tmp(17817) := x"ba60";
    tmp(17818) := x"b240";
    tmp(17819) := x"aa20";
    tmp(17820) := x"aa20";
    tmp(17821) := x"aa40";
    tmp(17822) := x"a220";
    tmp(17823) := x"a240";
    tmp(17824) := x"9200";
    tmp(17825) := x"89c0";
    tmp(17826) := x"6980";
    tmp(17827) := x"4100";
    tmp(17828) := x"28e0";
    tmp(17829) := x"18a0";
    tmp(17830) := x"1080";
    tmp(17831) := x"0860";
    tmp(17832) := x"0020";
    tmp(17833) := x"0000";
    tmp(17834) := x"0000";
    tmp(17835) := x"0000";
    tmp(17836) := x"0000";
    tmp(17837) := x"0000";
    tmp(17838) := x"0000";
    tmp(17839) := x"0000";
    tmp(17840) := x"0000";
    tmp(17841) := x"0000";
    tmp(17842) := x"0000";
    tmp(17843) := x"0000";
    tmp(17844) := x"0000";
    tmp(17845) := x"0000";
    tmp(17846) := x"0000";
    tmp(17847) := x"0000";
    tmp(17848) := x"0000";
    tmp(17849) := x"0000";
    tmp(17850) := x"0000";
    tmp(17851) := x"0000";
    tmp(17852) := x"0000";
    tmp(17853) := x"18a3";
    tmp(17854) := x"624a";
    tmp(17855) := x"5a09";
    tmp(17856) := x"59c8";
    tmp(17857) := x"724a";
    tmp(17858) := x"92cc";
    tmp(17859) := x"bbb1";
    tmp(17860) := x"c3f2";
    tmp(17861) := x"d475";
    tmp(17862) := x"e4f6";
    tmp(17863) := x"f558";
    tmp(17864) := x"fefe";
    tmp(17865) := x"fddb";
    tmp(17866) := x"fe9c";
    tmp(17867) := x"fede";
    tmp(17868) := x"e4f7";
    tmp(17869) := x"9aed";
    tmp(17870) := x"9aab";
    tmp(17871) := x"b36e";
    tmp(17872) := x"dc52";
    tmp(17873) := x"f536";
    tmp(17874) := x"fe3b";
    tmp(17875) := x"fefc";
    tmp(17876) := x"18a2";
    tmp(17877) := x"0020";
    tmp(17878) := x"0000";
    tmp(17879) := x"4185";
    tmp(17880) := x"ccf4";
    tmp(17881) := x"6269";
    tmp(17882) := x"0000";
    tmp(17883) := x"9bee";
    tmp(17884) := x"830d";
    tmp(17885) := x"1061";
    tmp(17886) := x"28e3";
    tmp(17887) := x"938f";
    tmp(17888) := x"9391";
    tmp(17889) := x"7b0f";
    tmp(17890) := x"7b0f";
    tmp(17891) := x"8bd1";
    tmp(17892) := x"3966";
    tmp(17893) := x"41e8";
    tmp(17894) := x"41c8";
    tmp(17895) := x"0821";
    tmp(17896) := x"5209";
    tmp(17897) := x"6b2c";
    tmp(17898) := x"0821";
    tmp(17899) := x"0000";
    tmp(17900) := x"20e3";
    tmp(17901) := x"736b";
    tmp(17902) := x"0881";
    tmp(17903) := x"0040";
    tmp(17904) := x"08a0";
    tmp(17905) := x"08c0";
    tmp(17906) := x"10e0";
    tmp(17907) := x"08c0";
    tmp(17908) := x"10e0";
    tmp(17909) := x"1120";
    tmp(17910) := x"1100";
    tmp(17911) := x"1960";
    tmp(17912) := x"19a0";
    tmp(17913) := x"2ac1";
    tmp(17914) := x"2241";
    tmp(17915) := x"19a0";
    tmp(17916) := x"08c0";
    tmp(17917) := x"08a0";
    tmp(17918) := x"08a0";
    tmp(17919) := x"08a0";
    tmp(17920) := x"08a0";
    tmp(17921) := x"08c0";
    tmp(17922) := x"10c0";
    tmp(17923) := x"10e0";
    tmp(17924) := x"18e1";
    tmp(17925) := x"1901";
    tmp(17926) := x"1901";
    tmp(17927) := x"2121";
    tmp(17928) := x"2141";
    tmp(17929) := x"2941";
    tmp(17930) := x"2961";
    tmp(17931) := x"3182";
    tmp(17932) := x"31a2";
    tmp(17933) := x"31a2";
    tmp(17934) := x"3181";
    tmp(17935) := x"2981";
    tmp(17936) := x"2981";
    tmp(17937) := x"2981";
    tmp(17938) := x"2981";
    tmp(17939) := x"2161";
    tmp(17940) := x"2161";
    tmp(17941) := x"2181";
    tmp(17942) := x"2161";
    tmp(17943) := x"2161";
    tmp(17944) := x"1961";
    tmp(17945) := x"1940";
    tmp(17946) := x"1940";
    tmp(17947) := x"1120";
    tmp(17948) := x"1100";
    tmp(17949) := x"10e0";
    tmp(17950) := x"08c0";
    tmp(17951) := x"08a0";
    tmp(17952) := x"0880";
    tmp(17953) := x"0860";
    tmp(17954) := x"0860";
    tmp(17955) := x"0860";
    tmp(17956) := x"0840";
    tmp(17957) := x"0000";
    tmp(17958) := x"0000";
    tmp(17959) := x"0000";
    tmp(17960) := x"0000";
    tmp(17961) := x"0000";
    tmp(17962) := x"0000";
    tmp(17963) := x"0000";
    tmp(17964) := x"0000";
    tmp(17965) := x"0000";
    tmp(17966) := x"0000";
    tmp(17967) := x"0000";
    tmp(17968) := x"0000";
    tmp(17969) := x"0000";
    tmp(17970) := x"0000";
    tmp(17971) := x"0000";
    tmp(17972) := x"0000";
    tmp(17973) := x"0000";
    tmp(17974) := x"0000";
    tmp(17975) := x"0000";
    tmp(17976) := x"0000";
    tmp(17977) := x"0000";
    tmp(17978) := x"0000";
    tmp(17979) := x"0000";
    tmp(17980) := x"0000";
    tmp(17981) := x"0000";
    tmp(17982) := x"0000";
    tmp(17983) := x"0000";
    tmp(17984) := x"0000";
    tmp(17985) := x"0000";
    tmp(17986) := x"0000";
    tmp(17987) := x"0000";
    tmp(17988) := x"0000";
    tmp(17989) := x"0000";
    tmp(17990) := x"0000";
    tmp(17991) := x"0000";
    tmp(17992) := x"0000";
    tmp(17993) := x"0000";
    tmp(17994) := x"0000";
    tmp(17995) := x"0000";
    tmp(17996) := x"0000";
    tmp(17997) := x"0840";
    tmp(17998) := x"0840";
    tmp(17999) := x"0840";
    tmp(18000) := x"1040";
    tmp(18001) := x"b260";
    tmp(18002) := x"a240";
    tmp(18003) := x"a240";
    tmp(18004) := x"a240";
    tmp(18005) := x"a260";
    tmp(18006) := x"aa60";
    tmp(18007) := x"b2a0";
    tmp(18008) := x"b2a0";
    tmp(18009) := x"baa0";
    tmp(18010) := x"baa0";
    tmp(18011) := x"c2c0";
    tmp(18012) := x"cb00";
    tmp(18013) := x"c2c0";
    tmp(18014) := x"cb20";
    tmp(18015) := x"db40";
    tmp(18016) := x"e340";
    tmp(18017) := x"db40";
    tmp(18018) := x"d320";
    tmp(18019) := x"d300";
    tmp(18020) := x"d2e0";
    tmp(18021) := x"e320";
    tmp(18022) := x"e300";
    tmp(18023) := x"e340";
    tmp(18024) := x"f3a0";
    tmp(18025) := x"f3a0";
    tmp(18026) := x"f380";
    tmp(18027) := x"eb80";
    tmp(18028) := x"fbc0";
    tmp(18029) := x"fbc0";
    tmp(18030) := x"fbe0";
    tmp(18031) := x"fc00";
    tmp(18032) := x"fc00";
    tmp(18033) := x"fc40";
    tmp(18034) := x"fc00";
    tmp(18035) := x"f400";
    tmp(18036) := x"e360";
    tmp(18037) := x"d2e0";
    tmp(18038) := x"cae0";
    tmp(18039) := x"cac0";
    tmp(18040) := x"ba80";
    tmp(18041) := x"b260";
    tmp(18042) := x"a240";
    tmp(18043) := x"aa40";
    tmp(18044) := x"a220";
    tmp(18045) := x"b260";
    tmp(18046) := x"b260";
    tmp(18047) := x"ba80";
    tmp(18048) := x"b280";
    tmp(18049) := x"b280";
    tmp(18050) := x"b260";
    tmp(18051) := x"aa40";
    tmp(18052) := x"aa20";
    tmp(18053) := x"aa40";
    tmp(18054) := x"b240";
    tmp(18055) := x"aa60";
    tmp(18056) := x"b260";
    tmp(18057) := x"ba80";
    tmp(18058) := x"b260";
    tmp(18059) := x"aa20";
    tmp(18060) := x"aa20";
    tmp(18061) := x"aa20";
    tmp(18062) := x"aa20";
    tmp(18063) := x"a220";
    tmp(18064) := x"9200";
    tmp(18065) := x"9200";
    tmp(18066) := x"7180";
    tmp(18067) := x"4920";
    tmp(18068) := x"28c0";
    tmp(18069) := x"1080";
    tmp(18070) := x"0860";
    tmp(18071) := x"0840";
    tmp(18072) := x"0020";
    tmp(18073) := x"0020";
    tmp(18074) := x"0000";
    tmp(18075) := x"0000";
    tmp(18076) := x"0000";
    tmp(18077) := x"0000";
    tmp(18078) := x"0000";
    tmp(18079) := x"0000";
    tmp(18080) := x"0000";
    tmp(18081) := x"0000";
    tmp(18082) := x"0000";
    tmp(18083) := x"0000";
    tmp(18084) := x"0000";
    tmp(18085) := x"0000";
    tmp(18086) := x"0000";
    tmp(18087) := x"0000";
    tmp(18088) := x"0000";
    tmp(18089) := x"0000";
    tmp(18090) := x"0000";
    tmp(18091) := x"0000";
    tmp(18092) := x"0000";
    tmp(18093) := x"1082";
    tmp(18094) := x"626a";
    tmp(18095) := x"59e8";
    tmp(18096) := x"6a29";
    tmp(18097) := x"7a6a";
    tmp(18098) := x"92cc";
    tmp(18099) := x"ab2e";
    tmp(18100) := x"bbb1";
    tmp(18101) := x"d494";
    tmp(18102) := x"dc94";
    tmp(18103) := x"ecf6";
    tmp(18104) := x"f6fd";
    tmp(18105) := x"f5b9";
    tmp(18106) := x"fefd";
    tmp(18107) := x"ff7f";
    tmp(18108) := x"ed78";
    tmp(18109) := x"b34f";
    tmp(18110) := x"a2cc";
    tmp(18111) := x"aaec";
    tmp(18112) := x"c36e";
    tmp(18113) := x"ecf4";
    tmp(18114) := x"fe5a";
    tmp(18115) := x"b410";
    tmp(18116) := x"0820";
    tmp(18117) := x"0000";
    tmp(18118) := x"0000";
    tmp(18119) := x"51e7";
    tmp(18120) := x"ed77";
    tmp(18121) := x"72cb";
    tmp(18122) := x"0820";
    tmp(18123) := x"d534";
    tmp(18124) := x"3945";
    tmp(18125) := x"0841";
    tmp(18126) := x"834d";
    tmp(18127) := x"9370";
    tmp(18128) := x"728d";
    tmp(18129) := x"28e5";
    tmp(18130) := x"20a3";
    tmp(18131) := x"3146";
    tmp(18132) := x"628c";
    tmp(18133) := x"5209";
    tmp(18134) := x"a432";
    tmp(18135) := x"49e8";
    tmp(18136) := x"0821";
    tmp(18137) := x"5aab";
    tmp(18138) := x"18a2";
    tmp(18139) := x"20e3";
    tmp(18140) := x"0841";
    tmp(18141) := x"2123";
    tmp(18142) := x"0860";
    tmp(18143) := x"0860";
    tmp(18144) := x"08a0";
    tmp(18145) := x"10e0";
    tmp(18146) := x"10e0";
    tmp(18147) := x"1100";
    tmp(18148) := x"1120";
    tmp(18149) := x"1960";
    tmp(18150) := x"1140";
    tmp(18151) := x"1980";
    tmp(18152) := x"2221";
    tmp(18153) := x"3342";
    tmp(18154) := x"2201";
    tmp(18155) := x"29c1";
    tmp(18156) := x"1941";
    tmp(18157) := x"1120";
    tmp(18158) := x"08e0";
    tmp(18159) := x"08a0";
    tmp(18160) := x"08a0";
    tmp(18161) := x"08a0";
    tmp(18162) := x"10c0";
    tmp(18163) := x"10e0";
    tmp(18164) := x"10e0";
    tmp(18165) := x"18e1";
    tmp(18166) := x"1901";
    tmp(18167) := x"1901";
    tmp(18168) := x"2101";
    tmp(18169) := x"2121";
    tmp(18170) := x"2941";
    tmp(18171) := x"2942";
    tmp(18172) := x"3162";
    tmp(18173) := x"3182";
    tmp(18174) := x"39a2";
    tmp(18175) := x"31a2";
    tmp(18176) := x"3181";
    tmp(18177) := x"2981";
    tmp(18178) := x"2981";
    tmp(18179) := x"2981";
    tmp(18180) := x"2981";
    tmp(18181) := x"2181";
    tmp(18182) := x"2181";
    tmp(18183) := x"2181";
    tmp(18184) := x"2181";
    tmp(18185) := x"2181";
    tmp(18186) := x"1961";
    tmp(18187) := x"1961";
    tmp(18188) := x"1940";
    tmp(18189) := x"1920";
    tmp(18190) := x"1100";
    tmp(18191) := x"10e0";
    tmp(18192) := x"08c0";
    tmp(18193) := x"08a0";
    tmp(18194) := x"0880";
    tmp(18195) := x"0860";
    tmp(18196) := x"0860";
    tmp(18197) := x"0000";
    tmp(18198) := x"0000";
    tmp(18199) := x"0000";
    tmp(18200) := x"0000";
    tmp(18201) := x"0000";
    tmp(18202) := x"0000";
    tmp(18203) := x"0000";
    tmp(18204) := x"0000";
    tmp(18205) := x"0000";
    tmp(18206) := x"0000";
    tmp(18207) := x"0000";
    tmp(18208) := x"0000";
    tmp(18209) := x"0000";
    tmp(18210) := x"0000";
    tmp(18211) := x"0000";
    tmp(18212) := x"0000";
    tmp(18213) := x"0000";
    tmp(18214) := x"0000";
    tmp(18215) := x"0000";
    tmp(18216) := x"0000";
    tmp(18217) := x"0000";
    tmp(18218) := x"0000";
    tmp(18219) := x"0000";
    tmp(18220) := x"0000";
    tmp(18221) := x"0000";
    tmp(18222) := x"0000";
    tmp(18223) := x"0000";
    tmp(18224) := x"0000";
    tmp(18225) := x"0000";
    tmp(18226) := x"0000";
    tmp(18227) := x"0000";
    tmp(18228) := x"0000";
    tmp(18229) := x"0000";
    tmp(18230) := x"0000";
    tmp(18231) := x"0000";
    tmp(18232) := x"0000";
    tmp(18233) := x"0000";
    tmp(18234) := x"0000";
    tmp(18235) := x"0000";
    tmp(18236) := x"0000";
    tmp(18237) := x"0840";
    tmp(18238) := x"0840";
    tmp(18239) := x"0840";
    tmp(18240) := x"1040";
    tmp(18241) := x"c2c0";
    tmp(18242) := x"b260";
    tmp(18243) := x"aa60";
    tmp(18244) := x"aa60";
    tmp(18245) := x"aa60";
    tmp(18246) := x"b280";
    tmp(18247) := x"ba80";
    tmp(18248) := x"baa0";
    tmp(18249) := x"baa0";
    tmp(18250) := x"bac0";
    tmp(18251) := x"c2c0";
    tmp(18252) := x"c2c0";
    tmp(18253) := x"c2c0";
    tmp(18254) := x"c2c0";
    tmp(18255) := x"d300";
    tmp(18256) := x"e340";
    tmp(18257) := x"db60";
    tmp(18258) := x"e360";
    tmp(18259) := x"e360";
    tmp(18260) := x"e340";
    tmp(18261) := x"eb80";
    tmp(18262) := x"e340";
    tmp(18263) := x"db20";
    tmp(18264) := x"eb60";
    tmp(18265) := x"f3a0";
    tmp(18266) := x"f380";
    tmp(18267) := x"f3a0";
    tmp(18268) := x"fc00";
    tmp(18269) := x"fc00";
    tmp(18270) := x"fbe0";
    tmp(18271) := x"fbe0";
    tmp(18272) := x"fbe0";
    tmp(18273) := x"fbe0";
    tmp(18274) := x"fb80";
    tmp(18275) := x"eb40";
    tmp(18276) := x"db00";
    tmp(18277) := x"cac0";
    tmp(18278) := x"d300";
    tmp(18279) := x"d300";
    tmp(18280) := x"cae0";
    tmp(18281) := x"baa0";
    tmp(18282) := x"aa40";
    tmp(18283) := x"aa40";
    tmp(18284) := x"b260";
    tmp(18285) := x"ba60";
    tmp(18286) := x"ba80";
    tmp(18287) := x"b260";
    tmp(18288) := x"ba60";
    tmp(18289) := x"aa60";
    tmp(18290) := x"a240";
    tmp(18291) := x"a220";
    tmp(18292) := x"a200";
    tmp(18293) := x"a200";
    tmp(18294) := x"aa40";
    tmp(18295) := x"b260";
    tmp(18296) := x"b280";
    tmp(18297) := x"ba80";
    tmp(18298) := x"ba80";
    tmp(18299) := x"a220";
    tmp(18300) := x"a200";
    tmp(18301) := x"a200";
    tmp(18302) := x"a200";
    tmp(18303) := x"a220";
    tmp(18304) := x"a220";
    tmp(18305) := x"9200";
    tmp(18306) := x"81c0";
    tmp(18307) := x"5960";
    tmp(18308) := x"30e0";
    tmp(18309) := x"1880";
    tmp(18310) := x"1080";
    tmp(18311) := x"0860";
    tmp(18312) := x"0840";
    tmp(18313) := x"0020";
    tmp(18314) := x"0000";
    tmp(18315) := x"0000";
    tmp(18316) := x"0000";
    tmp(18317) := x"0000";
    tmp(18318) := x"0000";
    tmp(18319) := x"0000";
    tmp(18320) := x"0000";
    tmp(18321) := x"0000";
    tmp(18322) := x"0000";
    tmp(18323) := x"0000";
    tmp(18324) := x"0000";
    tmp(18325) := x"0000";
    tmp(18326) := x"0000";
    tmp(18327) := x"0000";
    tmp(18328) := x"0000";
    tmp(18329) := x"0000";
    tmp(18330) := x"0000";
    tmp(18331) := x"0000";
    tmp(18332) := x"0000";
    tmp(18333) := x"0821";
    tmp(18334) := x"5229";
    tmp(18335) := x"5a09";
    tmp(18336) := x"6a29";
    tmp(18337) := x"7a4a";
    tmp(18338) := x"8a6b";
    tmp(18339) := x"ab4e";
    tmp(18340) := x"b34e";
    tmp(18341) := x"dc73";
    tmp(18342) := x"d472";
    tmp(18343) := x"f577";
    tmp(18344) := x"f579";
    tmp(18345) := x"f598";
    tmp(18346) := x"fedd";
    tmp(18347) := x"fe9b";
    tmp(18348) := x"ed57";
    tmp(18349) := x"c36f";
    tmp(18350) := x"c34e";
    tmp(18351) := x"c32e";
    tmp(18352) := x"cb8f";
    tmp(18353) := x"ecf4";
    tmp(18354) := x"fd97";
    tmp(18355) := x"932b";
    tmp(18356) := x"0820";
    tmp(18357) := x"0000";
    tmp(18358) := x"0020";
    tmp(18359) := x"934c";
    tmp(18360) := x"e597";
    tmp(18361) := x"3944";
    tmp(18362) := x"0841";
    tmp(18363) := x"a3f0";
    tmp(18364) := x"1882";
    tmp(18365) := x"18a2";
    tmp(18366) := x"9b8f";
    tmp(18367) := x"72ad";
    tmp(18368) := x"20c4";
    tmp(18369) := x"0820";
    tmp(18370) := x"0820";
    tmp(18371) := x"1062";
    tmp(18372) := x"18a3";
    tmp(18373) := x"520a";
    tmp(18374) := x"93b1";
    tmp(18375) := x"7aed";
    tmp(18376) := x"5248";
    tmp(18377) := x"0841";
    tmp(18378) := x"1082";
    tmp(18379) := x"5aaa";
    tmp(18380) := x"18c2";
    tmp(18381) := x"0020";
    tmp(18382) := x"0860";
    tmp(18383) := x"08a0";
    tmp(18384) := x"08c0";
    tmp(18385) := x"10e0";
    tmp(18386) := x"1100";
    tmp(18387) := x"1140";
    tmp(18388) := x"1140";
    tmp(18389) := x"1960";
    tmp(18390) := x"1960";
    tmp(18391) := x"1980";
    tmp(18392) := x"2a81";
    tmp(18393) := x"3342";
    tmp(18394) := x"3ac2";
    tmp(18395) := x"3a22";
    tmp(18396) := x"31c2";
    tmp(18397) := x"29a1";
    tmp(18398) := x"1961";
    tmp(18399) := x"1100";
    tmp(18400) := x"10e0";
    tmp(18401) := x"08c0";
    tmp(18402) := x"08c0";
    tmp(18403) := x"10c0";
    tmp(18404) := x"10e0";
    tmp(18405) := x"18e1";
    tmp(18406) := x"1901";
    tmp(18407) := x"1901";
    tmp(18408) := x"2101";
    tmp(18409) := x"2101";
    tmp(18410) := x"2121";
    tmp(18411) := x"2941";
    tmp(18412) := x"2942";
    tmp(18413) := x"3162";
    tmp(18414) := x"3982";
    tmp(18415) := x"39a2";
    tmp(18416) := x"39a2";
    tmp(18417) := x"31a2";
    tmp(18418) := x"3181";
    tmp(18419) := x"2981";
    tmp(18420) := x"29a1";
    tmp(18421) := x"29a1";
    tmp(18422) := x"29a1";
    tmp(18423) := x"29a1";
    tmp(18424) := x"29a1";
    tmp(18425) := x"29a1";
    tmp(18426) := x"29a1";
    tmp(18427) := x"21a1";
    tmp(18428) := x"2181";
    tmp(18429) := x"2161";
    tmp(18430) := x"1961";
    tmp(18431) := x"1921";
    tmp(18432) := x"1121";
    tmp(18433) := x"10e0";
    tmp(18434) := x"08a0";
    tmp(18435) := x"0880";
    tmp(18436) := x"0860";
    tmp(18437) := x"0000";
    tmp(18438) := x"0000";
    tmp(18439) := x"0000";
    tmp(18440) := x"0000";
    tmp(18441) := x"0000";
    tmp(18442) := x"0000";
    tmp(18443) := x"0000";
    tmp(18444) := x"0000";
    tmp(18445) := x"0000";
    tmp(18446) := x"0000";
    tmp(18447) := x"0000";
    tmp(18448) := x"0000";
    tmp(18449) := x"0000";
    tmp(18450) := x"0000";
    tmp(18451) := x"0000";
    tmp(18452) := x"0000";
    tmp(18453) := x"0000";
    tmp(18454) := x"0000";
    tmp(18455) := x"0000";
    tmp(18456) := x"0000";
    tmp(18457) := x"0000";
    tmp(18458) := x"0000";
    tmp(18459) := x"0000";
    tmp(18460) := x"0000";
    tmp(18461) := x"0000";
    tmp(18462) := x"0000";
    tmp(18463) := x"0000";
    tmp(18464) := x"0000";
    tmp(18465) := x"0000";
    tmp(18466) := x"0000";
    tmp(18467) := x"0000";
    tmp(18468) := x"0000";
    tmp(18469) := x"0000";
    tmp(18470) := x"0000";
    tmp(18471) := x"0000";
    tmp(18472) := x"0000";
    tmp(18473) := x"0000";
    tmp(18474) := x"0000";
    tmp(18475) := x"0000";
    tmp(18476) := x"0000";
    tmp(18477) := x"0840";
    tmp(18478) := x"0840";
    tmp(18479) := x"0840";
    tmp(18480) := x"1040";
    tmp(18481) := x"cac0";
    tmp(18482) := x"baa0";
    tmp(18483) := x"baa0";
    tmp(18484) := x"b280";
    tmp(18485) := x"bac0";
    tmp(18486) := x"baa0";
    tmp(18487) := x"ba80";
    tmp(18488) := x"c2a0";
    tmp(18489) := x"c2c0";
    tmp(18490) := x"c2e0";
    tmp(18491) := x"c2c0";
    tmp(18492) := x"c2e0";
    tmp(18493) := x"c2e0";
    tmp(18494) := x"c2c0";
    tmp(18495) := x"c2c0";
    tmp(18496) := x"cb00";
    tmp(18497) := x"db40";
    tmp(18498) := x"db40";
    tmp(18499) := x"db60";
    tmp(18500) := x"e360";
    tmp(18501) := x"eb80";
    tmp(18502) := x"eb80";
    tmp(18503) := x"e340";
    tmp(18504) := x"eb60";
    tmp(18505) := x"fbc0";
    tmp(18506) := x"fbc0";
    tmp(18507) := x"fbe0";
    tmp(18508) := x"fc00";
    tmp(18509) := x"fc20";
    tmp(18510) := x"fc00";
    tmp(18511) := x"fc20";
    tmp(18512) := x"fc40";
    tmp(18513) := x"fbe0";
    tmp(18514) := x"fb80";
    tmp(18515) := x"eb40";
    tmp(18516) := x"db00";
    tmp(18517) := x"d2e0";
    tmp(18518) := x"db20";
    tmp(18519) := x"db40";
    tmp(18520) := x"db20";
    tmp(18521) := x"cae0";
    tmp(18522) := x"b260";
    tmp(18523) := x"aa20";
    tmp(18524) := x"b260";
    tmp(18525) := x"b260";
    tmp(18526) := x"ba80";
    tmp(18527) := x"b280";
    tmp(18528) := x"b280";
    tmp(18529) := x"aa60";
    tmp(18530) := x"aa20";
    tmp(18531) := x"a220";
    tmp(18532) := x"a220";
    tmp(18533) := x"a220";
    tmp(18534) := x"aa40";
    tmp(18535) := x"b260";
    tmp(18536) := x"ba80";
    tmp(18537) := x"c2a0";
    tmp(18538) := x"ba60";
    tmp(18539) := x"aa20";
    tmp(18540) := x"a200";
    tmp(18541) := x"a200";
    tmp(18542) := x"9a00";
    tmp(18543) := x"a220";
    tmp(18544) := x"9a00";
    tmp(18545) := x"9a00";
    tmp(18546) := x"9a00";
    tmp(18547) := x"71a0";
    tmp(18548) := x"4100";
    tmp(18549) := x"20a0";
    tmp(18550) := x"1080";
    tmp(18551) := x"0860";
    tmp(18552) := x"0840";
    tmp(18553) := x"0020";
    tmp(18554) := x"0000";
    tmp(18555) := x"0000";
    tmp(18556) := x"0020";
    tmp(18557) := x"0000";
    tmp(18558) := x"0000";
    tmp(18559) := x"0000";
    tmp(18560) := x"0000";
    tmp(18561) := x"0000";
    tmp(18562) := x"0000";
    tmp(18563) := x"0000";
    tmp(18564) := x"0000";
    tmp(18565) := x"0000";
    tmp(18566) := x"0000";
    tmp(18567) := x"0000";
    tmp(18568) := x"0000";
    tmp(18569) := x"0000";
    tmp(18570) := x"0000";
    tmp(18571) := x"0000";
    tmp(18572) := x"0000";
    tmp(18573) := x"0000";
    tmp(18574) := x"18a3";
    tmp(18575) := x"624a";
    tmp(18576) := x"6a29";
    tmp(18577) := x"7a6a";
    tmp(18578) := x"8269";
    tmp(18579) := x"9acc";
    tmp(18580) := x"c3af";
    tmp(18581) := x"bb4d";
    tmp(18582) := x"dc72";
    tmp(18583) := x"ecf5";
    tmp(18584) := x"fd57";
    tmp(18585) := x"f4f5";
    tmp(18586) := x"fe39";
    tmp(18587) := x"fd98";
    tmp(18588) := x"ecf6";
    tmp(18589) := x"cb8f";
    tmp(18590) := x"d3d0";
    tmp(18591) := x"e431";
    tmp(18592) := x"dc10";
    tmp(18593) := x"f514";
    tmp(18594) := x"fd76";
    tmp(18595) := x"8b0b";
    tmp(18596) := x"0820";
    tmp(18597) := x"0000";
    tmp(18598) := x"0840";
    tmp(18599) := x"abce";
    tmp(18600) := x"dd15";
    tmp(18601) := x"1881";
    tmp(18602) := x"1882";
    tmp(18603) := x"7acb";
    tmp(18604) := x"18a2";
    tmp(18605) := x"5a08";
    tmp(18606) := x"7aed";
    tmp(18607) := x"2904";
    tmp(18608) := x"0841";
    tmp(18609) := x"18a2";
    tmp(18610) := x"41c6";
    tmp(18611) := x"41e6";
    tmp(18612) := x"2924";
    tmp(18613) := x"1882";
    tmp(18614) := x"41a7";
    tmp(18615) := x"9bd0";
    tmp(18616) := x"acb2";
    tmp(18617) := x"2924";
    tmp(18618) := x"18c2";
    tmp(18619) := x"18a2";
    tmp(18620) := x"10a2";
    tmp(18621) := x"0020";
    tmp(18622) := x"0880";
    tmp(18623) := x"08a0";
    tmp(18624) := x"08c0";
    tmp(18625) := x"10e0";
    tmp(18626) := x"1100";
    tmp(18627) := x"1140";
    tmp(18628) := x"1960";
    tmp(18629) := x"1140";
    tmp(18630) := x"1960";
    tmp(18631) := x"2200";
    tmp(18632) := x"2ae1";
    tmp(18633) := x"2a81";
    tmp(18634) := x"63c5";
    tmp(18635) := x"52c4";
    tmp(18636) := x"4a83";
    tmp(18637) := x"3a42";
    tmp(18638) := x"31e2";
    tmp(18639) := x"29a1";
    tmp(18640) := x"1961";
    tmp(18641) := x"1100";
    tmp(18642) := x"10e0";
    tmp(18643) := x"10c0";
    tmp(18644) := x"10c0";
    tmp(18645) := x"10e0";
    tmp(18646) := x"18e1";
    tmp(18647) := x"1901";
    tmp(18648) := x"1901";
    tmp(18649) := x"2101";
    tmp(18650) := x"2101";
    tmp(18651) := x"2921";
    tmp(18652) := x"2941";
    tmp(18653) := x"2942";
    tmp(18654) := x"3162";
    tmp(18655) := x"39a2";
    tmp(18656) := x"41c2";
    tmp(18657) := x"39a2";
    tmp(18658) := x"39a2";
    tmp(18659) := x"39a2";
    tmp(18660) := x"39c2";
    tmp(18661) := x"39e2";
    tmp(18662) := x"31e2";
    tmp(18663) := x"3a02";
    tmp(18664) := x"3202";
    tmp(18665) := x"3202";
    tmp(18666) := x"31e2";
    tmp(18667) := x"31e2";
    tmp(18668) := x"29e2";
    tmp(18669) := x"29a2";
    tmp(18670) := x"29a2";
    tmp(18671) := x"2181";
    tmp(18672) := x"2161";
    tmp(18673) := x"1941";
    tmp(18674) := x"1901";
    tmp(18675) := x"10e0";
    tmp(18676) := x"08a0";
    tmp(18677) := x"0000";
    tmp(18678) := x"0000";
    tmp(18679) := x"0000";
    tmp(18680) := x"0000";
    tmp(18681) := x"0000";
    tmp(18682) := x"0000";
    tmp(18683) := x"0000";
    tmp(18684) := x"0000";
    tmp(18685) := x"0000";
    tmp(18686) := x"0000";
    tmp(18687) := x"0000";
    tmp(18688) := x"0000";
    tmp(18689) := x"0000";
    tmp(18690) := x"0000";
    tmp(18691) := x"0000";
    tmp(18692) := x"0000";
    tmp(18693) := x"0000";
    tmp(18694) := x"0000";
    tmp(18695) := x"0000";
    tmp(18696) := x"0000";
    tmp(18697) := x"0000";
    tmp(18698) := x"0000";
    tmp(18699) := x"0000";
    tmp(18700) := x"0000";
    tmp(18701) := x"0000";
    tmp(18702) := x"0000";
    tmp(18703) := x"0000";
    tmp(18704) := x"0000";
    tmp(18705) := x"0000";
    tmp(18706) := x"0000";
    tmp(18707) := x"0000";
    tmp(18708) := x"0000";
    tmp(18709) := x"0000";
    tmp(18710) := x"0000";
    tmp(18711) := x"0000";
    tmp(18712) := x"0000";
    tmp(18713) := x"0000";
    tmp(18714) := x"0000";
    tmp(18715) := x"0000";
    tmp(18716) := x"0000";
    tmp(18717) := x"0840";
    tmp(18718) := x"0840";
    tmp(18719) := x"0840";
    tmp(18720) := x"1040";
    tmp(18721) := x"d300";
    tmp(18722) := x"c2c0";
    tmp(18723) := x"c2c0";
    tmp(18724) := x"c2c0";
    tmp(18725) := x"c2c0";
    tmp(18726) := x"c2a0";
    tmp(18727) := x"c2a0";
    tmp(18728) := x"cac0";
    tmp(18729) := x"cae0";
    tmp(18730) := x"c2e0";
    tmp(18731) := x"c2e0";
    tmp(18732) := x"c2c0";
    tmp(18733) := x"c2e0";
    tmp(18734) := x"c2c0";
    tmp(18735) := x"cac0";
    tmp(18736) := x"cae0";
    tmp(18737) := x"db20";
    tmp(18738) := x"db60";
    tmp(18739) := x"db60";
    tmp(18740) := x"e340";
    tmp(18741) := x"e340";
    tmp(18742) := x"e360";
    tmp(18743) := x"e360";
    tmp(18744) := x"eb80";
    tmp(18745) := x"fbc0";
    tmp(18746) := x"fbc0";
    tmp(18747) := x"fc00";
    tmp(18748) := x"fbe0";
    tmp(18749) := x"fc00";
    tmp(18750) := x"fc00";
    tmp(18751) := x"fc40";
    tmp(18752) := x"fc20";
    tmp(18753) := x"fbc0";
    tmp(18754) := x"eb60";
    tmp(18755) := x"e320";
    tmp(18756) := x"db00";
    tmp(18757) := x"d2e0";
    tmp(18758) := x"e340";
    tmp(18759) := x"eb40";
    tmp(18760) := x"e360";
    tmp(18761) := x"db40";
    tmp(18762) := x"c2a0";
    tmp(18763) := x"ba60";
    tmp(18764) := x"ba80";
    tmp(18765) := x"ba80";
    tmp(18766) := x"ba80";
    tmp(18767) := x"b260";
    tmp(18768) := x"ba80";
    tmp(18769) := x"b260";
    tmp(18770) := x"aa20";
    tmp(18771) := x"a220";
    tmp(18772) := x"aa40";
    tmp(18773) := x"aa40";
    tmp(18774) := x"b260";
    tmp(18775) := x"ba80";
    tmp(18776) := x"c2c0";
    tmp(18777) := x"c2c0";
    tmp(18778) := x"b260";
    tmp(18779) := x"aa40";
    tmp(18780) := x"a220";
    tmp(18781) := x"aa00";
    tmp(18782) := x"aa20";
    tmp(18783) := x"a220";
    tmp(18784) := x"9a20";
    tmp(18785) := x"a220";
    tmp(18786) := x"aa40";
    tmp(18787) := x"9200";
    tmp(18788) := x"5960";
    tmp(18789) := x"30e0";
    tmp(18790) := x"18a0";
    tmp(18791) := x"1060";
    tmp(18792) := x"0040";
    tmp(18793) := x"0020";
    tmp(18794) := x"0020";
    tmp(18795) := x"0020";
    tmp(18796) := x"0020";
    tmp(18797) := x"0020";
    tmp(18798) := x"0000";
    tmp(18799) := x"0000";
    tmp(18800) := x"0000";
    tmp(18801) := x"0000";
    tmp(18802) := x"0000";
    tmp(18803) := x"0000";
    tmp(18804) := x"0000";
    tmp(18805) := x"0000";
    tmp(18806) := x"0000";
    tmp(18807) := x"0000";
    tmp(18808) := x"0000";
    tmp(18809) := x"0000";
    tmp(18810) := x"0000";
    tmp(18811) := x"0000";
    tmp(18812) := x"0000";
    tmp(18813) := x"0000";
    tmp(18814) := x"0841";
    tmp(18815) := x"5a4a";
    tmp(18816) := x"6a6a";
    tmp(18817) := x"7229";
    tmp(18818) := x"7a49";
    tmp(18819) := x"928a";
    tmp(18820) := x"bb4d";
    tmp(18821) := x"bb4e";
    tmp(18822) := x"cb8f";
    tmp(18823) := x"ec92";
    tmp(18824) := x"f4f4";
    tmp(18825) := x"f4d5";
    tmp(18826) := x"fdb8";
    tmp(18827) := x"f4d5";
    tmp(18828) := x"e4d4";
    tmp(18829) := x"cbaf";
    tmp(18830) := x"e472";
    tmp(18831) := x"f556";
    tmp(18832) := x"f4d3";
    tmp(18833) := x"f596";
    tmp(18834) := x"fdf7";
    tmp(18835) := x"934b";
    tmp(18836) := x"0020";
    tmp(18837) := x"0000";
    tmp(18838) := x"4185";
    tmp(18839) := x"dd14";
    tmp(18840) := x"c472";
    tmp(18841) := x"0820";
    tmp(18842) := x"20a2";
    tmp(18843) := x"728a";
    tmp(18844) := x"20c3";
    tmp(18845) := x"6249";
    tmp(18846) := x"626a";
    tmp(18847) := x"1041";
    tmp(18848) := x"1061";
    tmp(18849) := x"41e5";
    tmp(18850) := x"41e6";
    tmp(18851) := x"3144";
    tmp(18852) := x"39a6";
    tmp(18853) := x"2945";
    tmp(18854) := x"0841";
    tmp(18855) := x"6a6a";
    tmp(18856) := x"936f";
    tmp(18857) := x"c5b6";
    tmp(18858) := x"41c6";
    tmp(18859) := x"0861";
    tmp(18860) := x"0020";
    tmp(18861) := x"0060";
    tmp(18862) := x"08a0";
    tmp(18863) := x"08c0";
    tmp(18864) := x"10e0";
    tmp(18865) := x"10e0";
    tmp(18866) := x"1100";
    tmp(18867) := x"1960";
    tmp(18868) := x"19a0";
    tmp(18869) := x"19a0";
    tmp(18870) := x"19e0";
    tmp(18871) := x"2261";
    tmp(18872) := x"2a61";
    tmp(18873) := x"42c3";
    tmp(18874) := x"8c88";
    tmp(18875) := x"7386";
    tmp(18876) := x"6325";
    tmp(18877) := x"52c4";
    tmp(18878) := x"4a83";
    tmp(18879) := x"3a22";
    tmp(18880) := x"31e2";
    tmp(18881) := x"2981";
    tmp(18882) := x"2161";
    tmp(18883) := x"1920";
    tmp(18884) := x"10e0";
    tmp(18885) := x"10e0";
    tmp(18886) := x"10e0";
    tmp(18887) := x"1901";
    tmp(18888) := x"1901";
    tmp(18889) := x"2101";
    tmp(18890) := x"2101";
    tmp(18891) := x"2101";
    tmp(18892) := x"2921";
    tmp(18893) := x"2941";
    tmp(18894) := x"3162";
    tmp(18895) := x"3982";
    tmp(18896) := x"41c3";
    tmp(18897) := x"4a03";
    tmp(18898) := x"4a03";
    tmp(18899) := x"4a03";
    tmp(18900) := x"4203";
    tmp(18901) := x"4a23";
    tmp(18902) := x"4223";
    tmp(18903) := x"4244";
    tmp(18904) := x"4244";
    tmp(18905) := x"4264";
    tmp(18906) := x"4243";
    tmp(18907) := x"4243";
    tmp(18908) := x"3a43";
    tmp(18909) := x"3a23";
    tmp(18910) := x"3203";
    tmp(18911) := x"31e3";
    tmp(18912) := x"29a2";
    tmp(18913) := x"29a2";
    tmp(18914) := x"2162";
    tmp(18915) := x"1941";
    tmp(18916) := x"1101";
    tmp(18917) := x"0000";
    tmp(18918) := x"0000";
    tmp(18919) := x"0000";
    tmp(18920) := x"0000";
    tmp(18921) := x"0000";
    tmp(18922) := x"0000";
    tmp(18923) := x"0000";
    tmp(18924) := x"0000";
    tmp(18925) := x"0000";
    tmp(18926) := x"0000";
    tmp(18927) := x"0000";
    tmp(18928) := x"0000";
    tmp(18929) := x"0000";
    tmp(18930) := x"0000";
    tmp(18931) := x"0000";
    tmp(18932) := x"0000";
    tmp(18933) := x"0000";
    tmp(18934) := x"0000";
    tmp(18935) := x"0000";
    tmp(18936) := x"0000";
    tmp(18937) := x"0000";
    tmp(18938) := x"0000";
    tmp(18939) := x"0000";
    tmp(18940) := x"0000";
    tmp(18941) := x"0000";
    tmp(18942) := x"0000";
    tmp(18943) := x"0000";
    tmp(18944) := x"0000";
    tmp(18945) := x"0000";
    tmp(18946) := x"0000";
    tmp(18947) := x"0000";
    tmp(18948) := x"0000";
    tmp(18949) := x"0000";
    tmp(18950) := x"0000";
    tmp(18951) := x"0000";
    tmp(18952) := x"0000";
    tmp(18953) := x"0000";
    tmp(18954) := x"0000";
    tmp(18955) := x"0000";
    tmp(18956) := x"0000";
    tmp(18957) := x"0840";
    tmp(18958) := x"0840";
    tmp(18959) := x"0840";
    tmp(18960) := x"1040";
    tmp(18961) := x"d320";
    tmp(18962) := x"c2c0";
    tmp(18963) := x"d2e0";
    tmp(18964) := x"d2e0";
    tmp(18965) := x"cac0";
    tmp(18966) := x"cac0";
    tmp(18967) := x"cac0";
    tmp(18968) := x"cac0";
    tmp(18969) := x"cac0";
    tmp(18970) := x"cae0";
    tmp(18971) := x"cae0";
    tmp(18972) := x"c2c0";
    tmp(18973) := x"baa0";
    tmp(18974) := x"baa0";
    tmp(18975) := x"cae0";
    tmp(18976) := x"d300";
    tmp(18977) := x"db40";
    tmp(18978) := x"db40";
    tmp(18979) := x"e360";
    tmp(18980) := x"e360";
    tmp(18981) := x"f380";
    tmp(18982) := x"f3a0";
    tmp(18983) := x"f3a0";
    tmp(18984) := x"f380";
    tmp(18985) := x"fba0";
    tmp(18986) := x"fba0";
    tmp(18987) := x"fbe0";
    tmp(18988) := x"fbe0";
    tmp(18989) := x"fc00";
    tmp(18990) := x"fbe0";
    tmp(18991) := x"fc00";
    tmp(18992) := x"fc40";
    tmp(18993) := x"fbe0";
    tmp(18994) := x"eb60";
    tmp(18995) := x"e300";
    tmp(18996) := x"dae0";
    tmp(18997) := x"db00";
    tmp(18998) := x"e340";
    tmp(18999) := x"eb60";
    tmp(19000) := x"e340";
    tmp(19001) := x"db20";
    tmp(19002) := x"cac0";
    tmp(19003) := x"caa0";
    tmp(19004) := x"c280";
    tmp(19005) := x"ba80";
    tmp(19006) := x"c2a0";
    tmp(19007) := x"ba80";
    tmp(19008) := x"baa0";
    tmp(19009) := x"b280";
    tmp(19010) := x"aa40";
    tmp(19011) := x"a220";
    tmp(19012) := x"aa20";
    tmp(19013) := x"b240";
    tmp(19014) := x"ba60";
    tmp(19015) := x"ba80";
    tmp(19016) := x"cac0";
    tmp(19017) := x"cae0";
    tmp(19018) := x"baa0";
    tmp(19019) := x"aa60";
    tmp(19020) := x"a220";
    tmp(19021) := x"9a00";
    tmp(19022) := x"a220";
    tmp(19023) := x"a200";
    tmp(19024) := x"a220";
    tmp(19025) := x"a220";
    tmp(19026) := x"a200";
    tmp(19027) := x"a240";
    tmp(19028) := x"89e0";
    tmp(19029) := x"4920";
    tmp(19030) := x"28c0";
    tmp(19031) := x"1080";
    tmp(19032) := x"0840";
    tmp(19033) := x"0020";
    tmp(19034) := x"0020";
    tmp(19035) := x"0020";
    tmp(19036) := x"0020";
    tmp(19037) := x"0020";
    tmp(19038) := x"0020";
    tmp(19039) := x"0000";
    tmp(19040) := x"0000";
    tmp(19041) := x"0000";
    tmp(19042) := x"0000";
    tmp(19043) := x"0000";
    tmp(19044) := x"0000";
    tmp(19045) := x"0000";
    tmp(19046) := x"0000";
    tmp(19047) := x"0000";
    tmp(19048) := x"0000";
    tmp(19049) := x"0000";
    tmp(19050) := x"0000";
    tmp(19051) := x"0000";
    tmp(19052) := x"0000";
    tmp(19053) := x"0000";
    tmp(19054) := x"0821";
    tmp(19055) := x"4187";
    tmp(19056) := x"7aed";
    tmp(19057) := x"7a8b";
    tmp(19058) := x"8aaa";
    tmp(19059) := x"9aab";
    tmp(19060) := x"a2ec";
    tmp(19061) := x"a2ec";
    tmp(19062) := x"b30c";
    tmp(19063) := x"e451";
    tmp(19064) := x"dc51";
    tmp(19065) := x"f4d4";
    tmp(19066) := x"ecd5";
    tmp(19067) := x"f516";
    tmp(19068) := x"e452";
    tmp(19069) := x"cb8f";
    tmp(19070) := x"dc31";
    tmp(19071) := x"fd56";
    tmp(19072) := x"fdf8";
    tmp(19073) := x"fe99";
    tmp(19074) := x"feb9";
    tmp(19075) := x"7b0a";
    tmp(19076) := x"0000";
    tmp(19077) := x"1041";
    tmp(19078) := x"ab8c";
    tmp(19079) := x"f5b7";
    tmp(19080) := x"b431";
    tmp(19081) := x"0820";
    tmp(19082) := x"1061";
    tmp(19083) := x"6a69";
    tmp(19084) := x"1861";
    tmp(19085) := x"49a7";
    tmp(19086) := x"51e8";
    tmp(19087) := x"0841";
    tmp(19088) := x"20c2";
    tmp(19089) := x"5226";
    tmp(19090) := x"20e3";
    tmp(19091) := x"0020";
    tmp(19092) := x"0841";
    tmp(19093) := x"31a6";
    tmp(19094) := x"18a2";
    tmp(19095) := x"1041";
    tmp(19096) := x"abf1";
    tmp(19097) := x"ddb7";
    tmp(19098) := x"944e";
    tmp(19099) := x"0840";
    tmp(19100) := x"0020";
    tmp(19101) := x"08a0";
    tmp(19102) := x"08c0";
    tmp(19103) := x"08c0";
    tmp(19104) := x"1100";
    tmp(19105) := x"1100";
    tmp(19106) := x"1120";
    tmp(19107) := x"1980";
    tmp(19108) := x"19a0";
    tmp(19109) := x"2260";
    tmp(19110) := x"1a00";
    tmp(19111) := x"2a81";
    tmp(19112) := x"21e1";
    tmp(19113) := x"9d49";
    tmp(19114) := x"9ca9";
    tmp(19115) := x"9469";
    tmp(19116) := x"83e7";
    tmp(19117) := x"7386";
    tmp(19118) := x"6345";
    tmp(19119) := x"5ae4";
    tmp(19120) := x"4a63";
    tmp(19121) := x"3a22";
    tmp(19122) := x"31e1";
    tmp(19123) := x"2981";
    tmp(19124) := x"2140";
    tmp(19125) := x"1900";
    tmp(19126) := x"10e0";
    tmp(19127) := x"10e0";
    tmp(19128) := x"1900";
    tmp(19129) := x"1901";
    tmp(19130) := x"2101";
    tmp(19131) := x"2101";
    tmp(19132) := x"2921";
    tmp(19133) := x"3141";
    tmp(19134) := x"3962";
    tmp(19135) := x"41a3";
    tmp(19136) := x"49e4";
    tmp(19137) := x"5a44";
    tmp(19138) := x"5a45";
    tmp(19139) := x"5a45";
    tmp(19140) := x"5245";
    tmp(19141) := x"5265";
    tmp(19142) := x"5265";
    tmp(19143) := x"5285";
    tmp(19144) := x"5285";
    tmp(19145) := x"5285";
    tmp(19146) := x"52a5";
    tmp(19147) := x"4a85";
    tmp(19148) := x"4a85";
    tmp(19149) := x"4265";
    tmp(19150) := x"4264";
    tmp(19151) := x"3a24";
    tmp(19152) := x"3204";
    tmp(19153) := x"31e4";
    tmp(19154) := x"31c3";
    tmp(19155) := x"29a3";
    tmp(19156) := x"2142";
    tmp(19157) := x"0000";
    tmp(19158) := x"0000";
    tmp(19159) := x"0000";
    tmp(19160) := x"0000";
    tmp(19161) := x"0000";
    tmp(19162) := x"0000";
    tmp(19163) := x"0000";
    tmp(19164) := x"0000";
    tmp(19165) := x"0000";
    tmp(19166) := x"0000";
    tmp(19167) := x"0000";
    tmp(19168) := x"0000";
    tmp(19169) := x"0000";
    tmp(19170) := x"0000";
    tmp(19171) := x"0000";
    tmp(19172) := x"0000";
    tmp(19173) := x"0000";
    tmp(19174) := x"0000";
    tmp(19175) := x"0000";
    tmp(19176) := x"0000";
    tmp(19177) := x"0000";
    tmp(19178) := x"0000";
    tmp(19179) := x"0000";
    tmp(19180) := x"0000";
    tmp(19181) := x"0000";
    tmp(19182) := x"0000";
    tmp(19183) := x"0000";
    tmp(19184) := x"0000";
    tmp(19185) := x"0000";
    tmp(19186) := x"0000";
    tmp(19187) := x"0000";
    tmp(19188) := x"0000";
    tmp(19189) := x"0000";
    tmp(19190) := x"0000";
    tmp(19191) := x"0000";
    tmp(19192) := x"0000";
    tmp(19193) := x"0000";
    tmp(19194) := x"0000";
    tmp(19195) := x"0000";
    tmp(19196) := x"0000";
    tmp(19197) := x"0840";
    tmp(19198) := x"0840";
    tmp(19199) := x"0840";
    tmp(19200) := x"1040";
    tmp(19201) := x"db00";
    tmp(19202) := x"cac0";
    tmp(19203) := x"db00";
    tmp(19204) := x"db20";
    tmp(19205) := x"e320";
    tmp(19206) := x"e320";
    tmp(19207) := x"db20";
    tmp(19208) := x"db00";
    tmp(19209) := x"dae0";
    tmp(19210) := x"db20";
    tmp(19211) := x"d300";
    tmp(19212) := x"cae0";
    tmp(19213) := x"c2c0";
    tmp(19214) := x"c2a0";
    tmp(19215) := x"cae0";
    tmp(19216) := x"d320";
    tmp(19217) := x"cb00";
    tmp(19218) := x"d320";
    tmp(19219) := x"db20";
    tmp(19220) := x"e360";
    tmp(19221) := x"eb80";
    tmp(19222) := x"f380";
    tmp(19223) := x"eb80";
    tmp(19224) := x"eb80";
    tmp(19225) := x"f3a0";
    tmp(19226) := x"fb80";
    tmp(19227) := x"fba0";
    tmp(19228) := x"fbe0";
    tmp(19229) := x"fbe0";
    tmp(19230) := x"fc00";
    tmp(19231) := x"fc20";
    tmp(19232) := x"fc00";
    tmp(19233) := x"fbc0";
    tmp(19234) := x"f360";
    tmp(19235) := x"eb40";
    tmp(19236) := x"db00";
    tmp(19237) := x"db00";
    tmp(19238) := x"e320";
    tmp(19239) := x"eb40";
    tmp(19240) := x"e340";
    tmp(19241) := x"e340";
    tmp(19242) := x"db20";
    tmp(19243) := x"d2c0";
    tmp(19244) := x"caa0";
    tmp(19245) := x"c280";
    tmp(19246) := x"c2a0";
    tmp(19247) := x"c2a0";
    tmp(19248) := x"ba80";
    tmp(19249) := x"aa60";
    tmp(19250) := x"aa40";
    tmp(19251) := x"aa40";
    tmp(19252) := x"b240";
    tmp(19253) := x"b260";
    tmp(19254) := x"ba60";
    tmp(19255) := x"ba80";
    tmp(19256) := x"cac0";
    tmp(19257) := x"cae0";
    tmp(19258) := x"bac0";
    tmp(19259) := x"b280";
    tmp(19260) := x"a220";
    tmp(19261) := x"91e0";
    tmp(19262) := x"9a00";
    tmp(19263) := x"a220";
    tmp(19264) := x"a220";
    tmp(19265) := x"a220";
    tmp(19266) := x"a200";
    tmp(19267) := x"aa20";
    tmp(19268) := x"9a20";
    tmp(19269) := x"71c0";
    tmp(19270) := x"4940";
    tmp(19271) := x"28c0";
    tmp(19272) := x"1060";
    tmp(19273) := x"0840";
    tmp(19274) := x"0020";
    tmp(19275) := x"0020";
    tmp(19276) := x"0020";
    tmp(19277) := x"0020";
    tmp(19278) := x"0020";
    tmp(19279) := x"0000";
    tmp(19280) := x"0000";
    tmp(19281) := x"0000";
    tmp(19282) := x"0000";
    tmp(19283) := x"0000";
    tmp(19284) := x"0000";
    tmp(19285) := x"0000";
    tmp(19286) := x"0000";
    tmp(19287) := x"0000";
    tmp(19288) := x"0000";
    tmp(19289) := x"0000";
    tmp(19290) := x"0000";
    tmp(19291) := x"0000";
    tmp(19292) := x"0000";
    tmp(19293) := x"0000";
    tmp(19294) := x"0020";
    tmp(19295) := x"18a3";
    tmp(19296) := x"6a8c";
    tmp(19297) := x"7aac";
    tmp(19298) := x"8aab";
    tmp(19299) := x"92aa";
    tmp(19300) := x"9aab";
    tmp(19301) := x"b34d";
    tmp(19302) := x"b30d";
    tmp(19303) := x"dbf0";
    tmp(19304) := x"bb2d";
    tmp(19305) := x"fcd4";
    tmp(19306) := x"dbaf";
    tmp(19307) := x"fcf6";
    tmp(19308) := x"d3d0";
    tmp(19309) := x"e3f0";
    tmp(19310) := x"ec31";
    tmp(19311) := x"f4d3";
    tmp(19312) := x"fdd6";
    tmp(19313) := x"fe78";
    tmp(19314) := x"fdf7";
    tmp(19315) := x"1081";
    tmp(19316) := x"0000";
    tmp(19317) := x"4164";
    tmp(19318) := x"dcb2";
    tmp(19319) := x"f535";
    tmp(19320) := x"a3ef";
    tmp(19321) := x"0000";
    tmp(19322) := x"20c2";
    tmp(19323) := x"6a69";
    tmp(19324) := x"1061";
    tmp(19325) := x"3924";
    tmp(19326) := x"51c7";
    tmp(19327) := x"0841";
    tmp(19328) := x"2903";
    tmp(19329) := x"5226";
    tmp(19330) := x"1081";
    tmp(19331) := x"0000";
    tmp(19332) := x"0000";
    tmp(19333) := x"18a3";
    tmp(19334) := x"2923";
    tmp(19335) := x"0820";
    tmp(19336) := x"938d";
    tmp(19337) := x"bc71";
    tmp(19338) := x"6b28";
    tmp(19339) := x"0020";
    tmp(19340) := x"0060";
    tmp(19341) := x"08a0";
    tmp(19342) := x"08e0";
    tmp(19343) := x"08e0";
    tmp(19344) := x"1120";
    tmp(19345) := x"1120";
    tmp(19346) := x"19a0";
    tmp(19347) := x"19e0";
    tmp(19348) := x"19c0";
    tmp(19349) := x"2281";
    tmp(19350) := x"22a1";
    tmp(19351) := x"2221";
    tmp(19352) := x"5ba4";
    tmp(19353) := x"c5ec";
    tmp(19354) := x"bd2b";
    tmp(19355) := x"b50b";
    tmp(19356) := x"a4ca";
    tmp(19357) := x"8c49";
    tmp(19358) := x"83e7";
    tmp(19359) := x"7366";
    tmp(19360) := x"6325";
    tmp(19361) := x"52c4";
    tmp(19362) := x"4a63";
    tmp(19363) := x"3a02";
    tmp(19364) := x"31c1";
    tmp(19365) := x"2981";
    tmp(19366) := x"1920";
    tmp(19367) := x"1100";
    tmp(19368) := x"10e0";
    tmp(19369) := x"1900";
    tmp(19370) := x"2121";
    tmp(19371) := x"2121";
    tmp(19372) := x"2941";
    tmp(19373) := x"3161";
    tmp(19374) := x"3982";
    tmp(19375) := x"41a3";
    tmp(19376) := x"5204";
    tmp(19377) := x"5a45";
    tmp(19378) := x"6286";
    tmp(19379) := x"6a86";
    tmp(19380) := x"62a6";
    tmp(19381) := x"6286";
    tmp(19382) := x"6286";
    tmp(19383) := x"5a86";
    tmp(19384) := x"5aa6";
    tmp(19385) := x"5aa6";
    tmp(19386) := x"52c6";
    tmp(19387) := x"52c6";
    tmp(19388) := x"52c6";
    tmp(19389) := x"52a6";
    tmp(19390) := x"4a85";
    tmp(19391) := x"4265";
    tmp(19392) := x"3a45";
    tmp(19393) := x"3a25";
    tmp(19394) := x"3a05";
    tmp(19395) := x"31e4";
    tmp(19396) := x"29a3";
    tmp(19397) := x"0000";
    tmp(19398) := x"0000";
    tmp(19399) := x"0000";
    tmp(19400) := x"0000";
    tmp(19401) := x"0000";
    tmp(19402) := x"0000";
    tmp(19403) := x"0000";
    tmp(19404) := x"0000";
    tmp(19405) := x"0000";
    tmp(19406) := x"0000";
    tmp(19407) := x"0000";
    tmp(19408) := x"0000";
    tmp(19409) := x"0000";
    tmp(19410) := x"0000";
    tmp(19411) := x"0000";
    tmp(19412) := x"0000";
    tmp(19413) := x"0000";
    tmp(19414) := x"0000";
    tmp(19415) := x"0000";
    tmp(19416) := x"0000";
    tmp(19417) := x"0000";
    tmp(19418) := x"0000";
    tmp(19419) := x"0000";
    tmp(19420) := x"0000";
    tmp(19421) := x"0000";
    tmp(19422) := x"0000";
    tmp(19423) := x"0000";
    tmp(19424) := x"0000";
    tmp(19425) := x"0000";
    tmp(19426) := x"0000";
    tmp(19427) := x"0000";
    tmp(19428) := x"0000";
    tmp(19429) := x"0000";
    tmp(19430) := x"0000";
    tmp(19431) := x"0000";
    tmp(19432) := x"0000";
    tmp(19433) := x"0000";
    tmp(19434) := x"0000";
    tmp(19435) := x"0000";
    tmp(19436) := x"0000";
    tmp(19437) := x"0840";
    tmp(19438) := x"0840";
    tmp(19439) := x"0840";
    tmp(19440) := x"1040";
    tmp(19441) := x"e320";
    tmp(19442) := x"dae0";
    tmp(19443) := x"d2e0";
    tmp(19444) := x"db00";
    tmp(19445) := x"eb00";
    tmp(19446) := x"eb20";
    tmp(19447) := x"f360";
    tmp(19448) := x"eb40";
    tmp(19449) := x"eb40";
    tmp(19450) := x"eb40";
    tmp(19451) := x"e340";
    tmp(19452) := x"db20";
    tmp(19453) := x"cac0";
    tmp(19454) := x"cac0";
    tmp(19455) := x"c2a0";
    tmp(19456) := x"cb00";
    tmp(19457) := x"cae0";
    tmp(19458) := x"cb00";
    tmp(19459) := x"db40";
    tmp(19460) := x"db40";
    tmp(19461) := x"e360";
    tmp(19462) := x"eb80";
    tmp(19463) := x"eb80";
    tmp(19464) := x"f3a0";
    tmp(19465) := x"f3c0";
    tmp(19466) := x"f380";
    tmp(19467) := x"eb60";
    tmp(19468) := x"fbe0";
    tmp(19469) := x"fbe0";
    tmp(19470) := x"fbe0";
    tmp(19471) := x"f3c0";
    tmp(19472) := x"eba0";
    tmp(19473) := x"eb60";
    tmp(19474) := x"eb40";
    tmp(19475) := x"eb40";
    tmp(19476) := x"db20";
    tmp(19477) := x"db00";
    tmp(19478) := x"e320";
    tmp(19479) := x"eb40";
    tmp(19480) := x"eb40";
    tmp(19481) := x"eb80";
    tmp(19482) := x"e340";
    tmp(19483) := x"cac0";
    tmp(19484) := x"cac0";
    tmp(19485) := x"cac0";
    tmp(19486) := x"cac0";
    tmp(19487) := x"c2c0";
    tmp(19488) := x"c2a0";
    tmp(19489) := x"b260";
    tmp(19490) := x"aa40";
    tmp(19491) := x"b240";
    tmp(19492) := x"b260";
    tmp(19493) := x"ba80";
    tmp(19494) := x"c2a0";
    tmp(19495) := x"c2a0";
    tmp(19496) := x"baa0";
    tmp(19497) := x"baa0";
    tmp(19498) := x"c2c0";
    tmp(19499) := x"b2a0";
    tmp(19500) := x"a240";
    tmp(19501) := x"9a20";
    tmp(19502) := x"aa40";
    tmp(19503) := x"a240";
    tmp(19504) := x"aa40";
    tmp(19505) := x"a240";
    tmp(19506) := x"a200";
    tmp(19507) := x"aa20";
    tmp(19508) := x"a220";
    tmp(19509) := x"8a00";
    tmp(19510) := x"6180";
    tmp(19511) := x"30e0";
    tmp(19512) := x"1880";
    tmp(19513) := x"0860";
    tmp(19514) := x"0840";
    tmp(19515) := x"0840";
    tmp(19516) := x"0840";
    tmp(19517) := x"0020";
    tmp(19518) := x"0020";
    tmp(19519) := x"0000";
    tmp(19520) := x"0000";
    tmp(19521) := x"0000";
    tmp(19522) := x"0000";
    tmp(19523) := x"0000";
    tmp(19524) := x"0020";
    tmp(19525) := x"0000";
    tmp(19526) := x"0000";
    tmp(19527) := x"0000";
    tmp(19528) := x"0000";
    tmp(19529) := x"0000";
    tmp(19530) := x"0000";
    tmp(19531) := x"0000";
    tmp(19532) := x"0000";
    tmp(19533) := x"0000";
    tmp(19534) := x"0000";
    tmp(19535) := x"0020";
    tmp(19536) := x"2904";
    tmp(19537) := x"8b6f";
    tmp(19538) := x"9b6e";
    tmp(19539) := x"92cb";
    tmp(19540) := x"8249";
    tmp(19541) := x"a2cb";
    tmp(19542) := x"aacb";
    tmp(19543) := x"d3af";
    tmp(19544) := x"d3cf";
    tmp(19545) := x"c32d";
    tmp(19546) := x"db8f";
    tmp(19547) := x"d3af";
    tmp(19548) := x"dbaf";
    tmp(19549) := x"cb4d";
    tmp(19550) := x"fc51";
    tmp(19551) := x"fcf2";
    tmp(19552) := x"fdf5";
    tmp(19553) := x"ff9d";
    tmp(19554) := x"3965";
    tmp(19555) := x"0000";
    tmp(19556) := x"0820";
    tmp(19557) := x"8aca";
    tmp(19558) := x"fe38";
    tmp(19559) := x"ed35";
    tmp(19560) := x"5207";
    tmp(19561) := x"0000";
    tmp(19562) := x"72ca";
    tmp(19563) := x"8b2c";
    tmp(19564) := x"1061";
    tmp(19565) := x"1861";
    tmp(19566) := x"6a6a";
    tmp(19567) := x"0841";
    tmp(19568) := x"1081";
    tmp(19569) := x"4a05";
    tmp(19570) := x"2923";
    tmp(19571) := x"0841";
    tmp(19572) := x"0840";
    tmp(19573) := x"18c2";
    tmp(19574) := x"3164";
    tmp(19575) := x"0820";
    tmp(19576) := x"72aa";
    tmp(19577) := x"93cc";
    tmp(19578) := x"10c1";
    tmp(19579) := x"0060";
    tmp(19580) := x"08a0";
    tmp(19581) := x"08a0";
    tmp(19582) := x"08e0";
    tmp(19583) := x"0900";
    tmp(19584) := x"1160";
    tmp(19585) := x"1120";
    tmp(19586) := x"1a00";
    tmp(19587) := x"19e0";
    tmp(19588) := x"1a00";
    tmp(19589) := x"19e1";
    tmp(19590) := x"2ae2";
    tmp(19591) := x"3282";
    tmp(19592) := x"ce8c";
    tmp(19593) := x"c56d";
    tmp(19594) := x"cd6d";
    tmp(19595) := x"c56d";
    tmp(19596) := x"bd4c";
    tmp(19597) := x"ad0b";
    tmp(19598) := x"a4ca";
    tmp(19599) := x"9449";
    tmp(19600) := x"7ba7";
    tmp(19601) := x"7366";
    tmp(19602) := x"6305";
    tmp(19603) := x"5283";
    tmp(19604) := x"4a63";
    tmp(19605) := x"3a02";
    tmp(19606) := x"31a1";
    tmp(19607) := x"2141";
    tmp(19608) := x"1900";
    tmp(19609) := x"18e0";
    tmp(19610) := x"1901";
    tmp(19611) := x"2121";
    tmp(19612) := x"2941";
    tmp(19613) := x"3182";
    tmp(19614) := x"39a2";
    tmp(19615) := x"41e3";
    tmp(19616) := x"4a04";
    tmp(19617) := x"5245";
    tmp(19618) := x"6286";
    tmp(19619) := x"6ac7";
    tmp(19620) := x"6ac7";
    tmp(19621) := x"6aa7";
    tmp(19622) := x"6aa7";
    tmp(19623) := x"6ac8";
    tmp(19624) := x"62e8";
    tmp(19625) := x"62e8";
    tmp(19626) := x"62e7";
    tmp(19627) := x"5ac7";
    tmp(19628) := x"5ae7";
    tmp(19629) := x"5ae7";
    tmp(19630) := x"5ae7";
    tmp(19631) := x"5286";
    tmp(19632) := x"4a86";
    tmp(19633) := x"4246";
    tmp(19634) := x"4226";
    tmp(19635) := x"3a25";
    tmp(19636) := x"3a05";
    tmp(19637) := x"0000";
    tmp(19638) := x"0000";
    tmp(19639) := x"0000";
    tmp(19640) := x"0000";
    tmp(19641) := x"0000";
    tmp(19642) := x"0000";
    tmp(19643) := x"0000";
    tmp(19644) := x"0000";
    tmp(19645) := x"0000";
    tmp(19646) := x"0000";
    tmp(19647) := x"0000";
    tmp(19648) := x"0000";
    tmp(19649) := x"0000";
    tmp(19650) := x"0000";
    tmp(19651) := x"0000";
    tmp(19652) := x"0000";
    tmp(19653) := x"0000";
    tmp(19654) := x"0000";
    tmp(19655) := x"0000";
    tmp(19656) := x"0000";
    tmp(19657) := x"0000";
    tmp(19658) := x"0000";
    tmp(19659) := x"0000";
    tmp(19660) := x"0000";
    tmp(19661) := x"0000";
    tmp(19662) := x"0000";
    tmp(19663) := x"0000";
    tmp(19664) := x"0000";
    tmp(19665) := x"0000";
    tmp(19666) := x"0000";
    tmp(19667) := x"0000";
    tmp(19668) := x"0000";
    tmp(19669) := x"0000";
    tmp(19670) := x"0000";
    tmp(19671) := x"0000";
    tmp(19672) := x"0000";
    tmp(19673) := x"0000";
    tmp(19674) := x"0000";
    tmp(19675) := x"0000";
    tmp(19676) := x"0000";
    tmp(19677) := x"0840";
    tmp(19678) := x"0840";
    tmp(19679) := x"0840";
    tmp(19680) := x"1840";
    tmp(19681) := x"eb20";
    tmp(19682) := x"db00";
    tmp(19683) := x"db00";
    tmp(19684) := x"e300";
    tmp(19685) := x"e300";
    tmp(19686) := x"f340";
    tmp(19687) := x"f340";
    tmp(19688) := x"f340";
    tmp(19689) := x"fb60";
    tmp(19690) := x"fba0";
    tmp(19691) := x"fbc0";
    tmp(19692) := x"eb60";
    tmp(19693) := x"d2e0";
    tmp(19694) := x"cac0";
    tmp(19695) := x"cac0";
    tmp(19696) := x"cae0";
    tmp(19697) := x"cae0";
    tmp(19698) := x"d320";
    tmp(19699) := x"d320";
    tmp(19700) := x"d340";
    tmp(19701) := x"db40";
    tmp(19702) := x"e340";
    tmp(19703) := x"eb80";
    tmp(19704) := x"eb80";
    tmp(19705) := x"db40";
    tmp(19706) := x"eb40";
    tmp(19707) := x"eb60";
    tmp(19708) := x"eb60";
    tmp(19709) := x"f3c0";
    tmp(19710) := x"f3a0";
    tmp(19711) := x"fbc0";
    tmp(19712) := x"eb80";
    tmp(19713) := x"eb60";
    tmp(19714) := x"eb40";
    tmp(19715) := x"f360";
    tmp(19716) := x"e320";
    tmp(19717) := x"e300";
    tmp(19718) := x"eb20";
    tmp(19719) := x"eb20";
    tmp(19720) := x"eb40";
    tmp(19721) := x"eb40";
    tmp(19722) := x"eb60";
    tmp(19723) := x"db20";
    tmp(19724) := x"db00";
    tmp(19725) := x"d300";
    tmp(19726) := x"cac0";
    tmp(19727) := x"ba80";
    tmp(19728) := x"ba80";
    tmp(19729) := x"b240";
    tmp(19730) := x"aa40";
    tmp(19731) := x"aa40";
    tmp(19732) := x"b260";
    tmp(19733) := x"ba80";
    tmp(19734) := x"ba60";
    tmp(19735) := x"c2a0";
    tmp(19736) := x"cae0";
    tmp(19737) := x"c2e0";
    tmp(19738) := x"cb00";
    tmp(19739) := x"b280";
    tmp(19740) := x"a220";
    tmp(19741) := x"a240";
    tmp(19742) := x"aa20";
    tmp(19743) := x"aa40";
    tmp(19744) := x"aa40";
    tmp(19745) := x"aa40";
    tmp(19746) := x"a200";
    tmp(19747) := x"a220";
    tmp(19748) := x"a220";
    tmp(19749) := x"81c0";
    tmp(19750) := x"6160";
    tmp(19751) := x"4100";
    tmp(19752) := x"20c0";
    tmp(19753) := x"1080";
    tmp(19754) := x"0860";
    tmp(19755) := x"0860";
    tmp(19756) := x"0020";
    tmp(19757) := x"0020";
    tmp(19758) := x"0020";
    tmp(19759) := x"0020";
    tmp(19760) := x"0000";
    tmp(19761) := x"0000";
    tmp(19762) := x"0000";
    tmp(19763) := x"0000";
    tmp(19764) := x"0020";
    tmp(19765) := x"0000";
    tmp(19766) := x"0000";
    tmp(19767) := x"0000";
    tmp(19768) := x"0000";
    tmp(19769) := x"0000";
    tmp(19770) := x"0000";
    tmp(19771) := x"0000";
    tmp(19772) := x"0000";
    tmp(19773) := x"0000";
    tmp(19774) := x"0000";
    tmp(19775) := x"0000";
    tmp(19776) := x"0020";
    tmp(19777) := x"1082";
    tmp(19778) := x"5a08";
    tmp(19779) := x"a38f";
    tmp(19780) := x"7a49";
    tmp(19781) := x"8a69";
    tmp(19782) := x"b32c";
    tmp(19783) := x"aacb";
    tmp(19784) := x"cb6e";
    tmp(19785) := x"c34d";
    tmp(19786) := x"cb6e";
    tmp(19787) := x"bb0c";
    tmp(19788) := x"d36d";
    tmp(19789) := x"db8e";
    tmp(19790) := x"f4b1";
    tmp(19791) := x"fdb4";
    tmp(19792) := x"fed9";
    tmp(19793) := x"8b8d";
    tmp(19794) := x"0820";
    tmp(19795) := x"0000";
    tmp(19796) := x"20c2";
    tmp(19797) := x"c430";
    tmp(19798) := x"fd95";
    tmp(19799) := x"dd14";
    tmp(19800) := x"0820";
    tmp(19801) := x"1041";
    tmp(19802) := x"d4f3";
    tmp(19803) := x"b451";
    tmp(19804) := x"2903";
    tmp(19805) := x"0841";
    tmp(19806) := x"6a69";
    tmp(19807) := x"28e3";
    tmp(19808) := x"0820";
    tmp(19809) := x"2903";
    tmp(19810) := x"5246";
    tmp(19811) := x"3984";
    tmp(19812) := x"3143";
    tmp(19813) := x"39a5";
    tmp(19814) := x"2943";
    tmp(19815) := x"0820";
    tmp(19816) := x"6a68";
    tmp(19817) := x"5265";
    tmp(19818) := x"0860";
    tmp(19819) := x"0880";
    tmp(19820) := x"08e0";
    tmp(19821) := x"08e0";
    tmp(19822) := x"0900";
    tmp(19823) := x"1140";
    tmp(19824) := x"1180";
    tmp(19825) := x"1180";
    tmp(19826) := x"19e0";
    tmp(19827) := x"1a01";
    tmp(19828) := x"1a22";
    tmp(19829) := x"1a42";
    tmp(19830) := x"2201";
    tmp(19831) := x"7c87";
    tmp(19832) := x"bd2c";
    tmp(19833) := x"c56d";
    tmp(19834) := x"cdae";
    tmp(19835) := x"cdae";
    tmp(19836) := x"cdae";
    tmp(19837) := x"cd8d";
    tmp(19838) := x"bd4c";
    tmp(19839) := x"accb";
    tmp(19840) := x"9c8a";
    tmp(19841) := x"9428";
    tmp(19842) := x"7b87";
    tmp(19843) := x"6b25";
    tmp(19844) := x"62e4";
    tmp(19845) := x"5283";
    tmp(19846) := x"4242";
    tmp(19847) := x"31e1";
    tmp(19848) := x"2981";
    tmp(19849) := x"1920";
    tmp(19850) := x"1900";
    tmp(19851) := x"2121";
    tmp(19852) := x"2961";
    tmp(19853) := x"3182";
    tmp(19854) := x"39c2";
    tmp(19855) := x"41e4";
    tmp(19856) := x"4a04";
    tmp(19857) := x"5225";
    tmp(19858) := x"5a66";
    tmp(19859) := x"6aa7";
    tmp(19860) := x"72c7";
    tmp(19861) := x"6ac8";
    tmp(19862) := x"6ac8";
    tmp(19863) := x"6ac8";
    tmp(19864) := x"6ae9";
    tmp(19865) := x"6ae9";
    tmp(19866) := x"6b09";
    tmp(19867) := x"6ae9";
    tmp(19868) := x"6b09";
    tmp(19869) := x"6308";
    tmp(19870) := x"6308";
    tmp(19871) := x"5b08";
    tmp(19872) := x"52a7";
    tmp(19873) := x"52a7";
    tmp(19874) := x"4a87";
    tmp(19875) := x"4247";
    tmp(19876) := x"4246";
    tmp(19877) := x"0000";
    tmp(19878) := x"0000";
    tmp(19879) := x"0000";
    tmp(19880) := x"0000";
    tmp(19881) := x"0000";
    tmp(19882) := x"0000";
    tmp(19883) := x"0000";
    tmp(19884) := x"0000";
    tmp(19885) := x"0000";
    tmp(19886) := x"0000";
    tmp(19887) := x"0000";
    tmp(19888) := x"0000";
    tmp(19889) := x"0000";
    tmp(19890) := x"0000";
    tmp(19891) := x"0000";
    tmp(19892) := x"0000";
    tmp(19893) := x"0000";
    tmp(19894) := x"0000";
    tmp(19895) := x"0000";
    tmp(19896) := x"0000";
    tmp(19897) := x"0000";
    tmp(19898) := x"0000";
    tmp(19899) := x"0000";
    tmp(19900) := x"0000";
    tmp(19901) := x"0000";
    tmp(19902) := x"0000";
    tmp(19903) := x"0000";
    tmp(19904) := x"0000";
    tmp(19905) := x"0000";
    tmp(19906) := x"0000";
    tmp(19907) := x"0000";
    tmp(19908) := x"0000";
    tmp(19909) := x"0000";
    tmp(19910) := x"0000";
    tmp(19911) := x"0000";
    tmp(19912) := x"0000";
    tmp(19913) := x"0000";
    tmp(19914) := x"0000";
    tmp(19915) := x"0000";
    tmp(19916) := x"0000";
    tmp(19917) := x"0840";
    tmp(19918) := x"0840";
    tmp(19919) := x"0840";
    tmp(19920) := x"1040";
    tmp(19921) := x"f340";
    tmp(19922) := x"e320";
    tmp(19923) := x"e300";
    tmp(19924) := x"e300";
    tmp(19925) := x"eb00";
    tmp(19926) := x"eb20";
    tmp(19927) := x"f320";
    tmp(19928) := x"f340";
    tmp(19929) := x"fb40";
    tmp(19930) := x"fb60";
    tmp(19931) := x"f360";
    tmp(19932) := x"fba0";
    tmp(19933) := x"f3a0";
    tmp(19934) := x"d2e0";
    tmp(19935) := x"d2c0";
    tmp(19936) := x"d300";
    tmp(19937) := x"cae0";
    tmp(19938) := x"cb20";
    tmp(19939) := x"d320";
    tmp(19940) := x"db20";
    tmp(19941) := x"db40";
    tmp(19942) := x"db20";
    tmp(19943) := x"e340";
    tmp(19944) := x"eb80";
    tmp(19945) := x"db20";
    tmp(19946) := x"e340";
    tmp(19947) := x"e360";
    tmp(19948) := x"eb80";
    tmp(19949) := x"eb80";
    tmp(19950) := x"eba0";
    tmp(19951) := x"f3a0";
    tmp(19952) := x"fba0";
    tmp(19953) := x"eb60";
    tmp(19954) := x"eb60";
    tmp(19955) := x"eb80";
    tmp(19956) := x"e340";
    tmp(19957) := x"e300";
    tmp(19958) := x"eb20";
    tmp(19959) := x"eb20";
    tmp(19960) := x"eb40";
    tmp(19961) := x"eb40";
    tmp(19962) := x"f360";
    tmp(19963) := x"fb80";
    tmp(19964) := x"f360";
    tmp(19965) := x"e320";
    tmp(19966) := x"db00";
    tmp(19967) := x"cac0";
    tmp(19968) := x"caa0";
    tmp(19969) := x"ba60";
    tmp(19970) := x"b240";
    tmp(19971) := x"b240";
    tmp(19972) := x"ba60";
    tmp(19973) := x"c280";
    tmp(19974) := x"c2a0";
    tmp(19975) := x"c2c0";
    tmp(19976) := x"cb00";
    tmp(19977) := x"cb00";
    tmp(19978) := x"cb00";
    tmp(19979) := x"baa0";
    tmp(19980) := x"aa60";
    tmp(19981) := x"b260";
    tmp(19982) := x"a200";
    tmp(19983) := x"aa20";
    tmp(19984) := x"aa40";
    tmp(19985) := x"aa40";
    tmp(19986) := x"aa20";
    tmp(19987) := x"aa40";
    tmp(19988) := x"aa40";
    tmp(19989) := x"9a00";
    tmp(19990) := x"81c0";
    tmp(19991) := x"6160";
    tmp(19992) := x"3900";
    tmp(19993) := x"18a0";
    tmp(19994) := x"0860";
    tmp(19995) := x"0840";
    tmp(19996) := x"0860";
    tmp(19997) := x"0840";
    tmp(19998) := x"0020";
    tmp(19999) := x"0020";
    tmp(20000) := x"0000";
    tmp(20001) := x"0000";
    tmp(20002) := x"0000";
    tmp(20003) := x"0020";
    tmp(20004) := x"0000";
    tmp(20005) := x"0000";
    tmp(20006) := x"0000";
    tmp(20007) := x"0000";
    tmp(20008) := x"0000";
    tmp(20009) := x"0000";
    tmp(20010) := x"0000";
    tmp(20011) := x"0000";
    tmp(20012) := x"0000";
    tmp(20013) := x"0000";
    tmp(20014) := x"0000";
    tmp(20015) := x"0000";
    tmp(20016) := x"0000";
    tmp(20017) := x"0000";
    tmp(20018) := x"0841";
    tmp(20019) := x"624a";
    tmp(20020) := x"9b8e";
    tmp(20021) := x"8aeb";
    tmp(20022) := x"a30c";
    tmp(20023) := x"bb6d";
    tmp(20024) := x"aaeb";
    tmp(20025) := x"b32c";
    tmp(20026) := x"9a8a";
    tmp(20027) := x"bb0c";
    tmp(20028) := x"baeb";
    tmp(20029) := x"ebef";
    tmp(20030) := x"dc0f";
    tmp(20031) := x"fed8";
    tmp(20032) := x"b4d2";
    tmp(20033) := x"0841";
    tmp(20034) := x"0000";
    tmp(20035) := x"1081";
    tmp(20036) := x"b3ed";
    tmp(20037) := x"f553";
    tmp(20038) := x"fe99";
    tmp(20039) := x"1882";
    tmp(20040) := x"0000";
    tmp(20041) := x"6227";
    tmp(20042) := x"d4d3";
    tmp(20043) := x"bc93";
    tmp(20044) := x"5a49";
    tmp(20045) := x"0820";
    tmp(20046) := x"20a2";
    tmp(20047) := x"728a";
    tmp(20048) := x"20c3";
    tmp(20049) := x"0820";
    tmp(20050) := x"1081";
    tmp(20051) := x"3143";
    tmp(20052) := x"39a4";
    tmp(20053) := x"20c2";
    tmp(20054) := x"0020";
    tmp(20055) := x"18a2";
    tmp(20056) := x"6a88";
    tmp(20057) := x"1901";
    tmp(20058) := x"0860";
    tmp(20059) := x"08a0";
    tmp(20060) := x"08c0";
    tmp(20061) := x"0900";
    tmp(20062) := x"1120";
    tmp(20063) := x"1180";
    tmp(20064) := x"11a0";
    tmp(20065) := x"19c0";
    tmp(20066) := x"19e0";
    tmp(20067) := x"19e1";
    tmp(20068) := x"22a4";
    tmp(20069) := x"22c4";
    tmp(20070) := x"4303";
    tmp(20071) := x"ad2a";
    tmp(20072) := x"b4cb";
    tmp(20073) := x"c52d";
    tmp(20074) := x"cdae";
    tmp(20075) := x"d5cf";
    tmp(20076) := x"ddef";
    tmp(20077) := x"ddee";
    tmp(20078) := x"ddee";
    tmp(20079) := x"cd6d";
    tmp(20080) := x"b52b";
    tmp(20081) := x"acea";
    tmp(20082) := x"9449";
    tmp(20083) := x"8c08";
    tmp(20084) := x"7b66";
    tmp(20085) := x"6b25";
    tmp(20086) := x"5aa4";
    tmp(20087) := x"4a63";
    tmp(20088) := x"3a02";
    tmp(20089) := x"29a1";
    tmp(20090) := x"2141";
    tmp(20091) := x"2121";
    tmp(20092) := x"2141";
    tmp(20093) := x"2982";
    tmp(20094) := x"39c3";
    tmp(20095) := x"4204";
    tmp(20096) := x"4a04";
    tmp(20097) := x"5245";
    tmp(20098) := x"5a66";
    tmp(20099) := x"62a7";
    tmp(20100) := x"72e8";
    tmp(20101) := x"72e9";
    tmp(20102) := x"72c9";
    tmp(20103) := x"7b0a";
    tmp(20104) := x"7b2a";
    tmp(20105) := x"730a";
    tmp(20106) := x"732a";
    tmp(20107) := x"732a";
    tmp(20108) := x"732a";
    tmp(20109) := x"734a";
    tmp(20110) := x"6b4a";
    tmp(20111) := x"6b29";
    tmp(20112) := x"6308";
    tmp(20113) := x"52c8";
    tmp(20114) := x"52c8";
    tmp(20115) := x"4a88";
    tmp(20116) := x"4268";
    tmp(20117) := x"0000";
    tmp(20118) := x"0000";
    tmp(20119) := x"0000";
    tmp(20120) := x"0000";
    tmp(20121) := x"0000";
    tmp(20122) := x"0000";
    tmp(20123) := x"0000";
    tmp(20124) := x"0000";
    tmp(20125) := x"0000";
    tmp(20126) := x"0000";
    tmp(20127) := x"0000";
    tmp(20128) := x"0000";
    tmp(20129) := x"0000";
    tmp(20130) := x"0000";
    tmp(20131) := x"0000";
    tmp(20132) := x"0000";
    tmp(20133) := x"0000";
    tmp(20134) := x"0000";
    tmp(20135) := x"0000";
    tmp(20136) := x"0000";
    tmp(20137) := x"0000";
    tmp(20138) := x"0000";
    tmp(20139) := x"0000";
    tmp(20140) := x"0000";
    tmp(20141) := x"0000";
    tmp(20142) := x"0000";
    tmp(20143) := x"0000";
    tmp(20144) := x"0000";
    tmp(20145) := x"0000";
    tmp(20146) := x"0000";
    tmp(20147) := x"0000";
    tmp(20148) := x"0000";
    tmp(20149) := x"0000";
    tmp(20150) := x"0000";
    tmp(20151) := x"0000";
    tmp(20152) := x"0000";
    tmp(20153) := x"0000";
    tmp(20154) := x"0000";
    tmp(20155) := x"0000";
    tmp(20156) := x"0000";
    tmp(20157) := x"0840";
    tmp(20158) := x"0840";
    tmp(20159) := x"0840";
    tmp(20160) := x"1040";
    tmp(20161) := x"eb40";
    tmp(20162) := x"dae0";
    tmp(20163) := x"eb40";
    tmp(20164) := x"eb40";
    tmp(20165) := x"f340";
    tmp(20166) := x"eb20";
    tmp(20167) := x"f320";
    tmp(20168) := x"f340";
    tmp(20169) := x"f360";
    tmp(20170) := x"fb60";
    tmp(20171) := x"f360";
    tmp(20172) := x"f360";
    tmp(20173) := x"fb80";
    tmp(20174) := x"e300";
    tmp(20175) := x"e320";
    tmp(20176) := x"db20";
    tmp(20177) := x"d300";
    tmp(20178) := x"cae0";
    tmp(20179) := x"d300";
    tmp(20180) := x"e340";
    tmp(20181) := x"e340";
    tmp(20182) := x"db40";
    tmp(20183) := x"db40";
    tmp(20184) := x"db20";
    tmp(20185) := x"db00";
    tmp(20186) := x"d300";
    tmp(20187) := x"db20";
    tmp(20188) := x"eb80";
    tmp(20189) := x"f380";
    tmp(20190) := x"eb80";
    tmp(20191) := x"f3e0";
    tmp(20192) := x"f3a0";
    tmp(20193) := x"f360";
    tmp(20194) := x"eb40";
    tmp(20195) := x"f360";
    tmp(20196) := x"f360";
    tmp(20197) := x"f340";
    tmp(20198) := x"eb40";
    tmp(20199) := x"eb40";
    tmp(20200) := x"eb40";
    tmp(20201) := x"eb60";
    tmp(20202) := x"f380";
    tmp(20203) := x"fb80";
    tmp(20204) := x"fb80";
    tmp(20205) := x"fbc0";
    tmp(20206) := x"f360";
    tmp(20207) := x"db00";
    tmp(20208) := x"c2a0";
    tmp(20209) := x"b240";
    tmp(20210) := x"aa20";
    tmp(20211) := x"b240";
    tmp(20212) := x"c280";
    tmp(20213) := x"c280";
    tmp(20214) := x"c280";
    tmp(20215) := x"d2c0";
    tmp(20216) := x"db00";
    tmp(20217) := x"db20";
    tmp(20218) := x"cb00";
    tmp(20219) := x"c2e0";
    tmp(20220) := x"b260";
    tmp(20221) := x"a220";
    tmp(20222) := x"aa20";
    tmp(20223) := x"b260";
    tmp(20224) := x"b240";
    tmp(20225) := x"b260";
    tmp(20226) := x"b260";
    tmp(20227) := x"aa40";
    tmp(20228) := x"a220";
    tmp(20229) := x"a240";
    tmp(20230) := x"79a0";
    tmp(20231) := x"5940";
    tmp(20232) := x"4100";
    tmp(20233) := x"28c0";
    tmp(20234) := x"18a0";
    tmp(20235) := x"1080";
    tmp(20236) := x"1060";
    tmp(20237) := x"0860";
    tmp(20238) := x"0840";
    tmp(20239) := x"0840";
    tmp(20240) := x"0020";
    tmp(20241) := x"0000";
    tmp(20242) := x"0000";
    tmp(20243) := x"0000";
    tmp(20244) := x"0000";
    tmp(20245) := x"0000";
    tmp(20246) := x"0020";
    tmp(20247) := x"0020";
    tmp(20248) := x"0020";
    tmp(20249) := x"0000";
    tmp(20250) := x"0000";
    tmp(20251) := x"0000";
    tmp(20252) := x"0000";
    tmp(20253) := x"0000";
    tmp(20254) := x"0000";
    tmp(20255) := x"0000";
    tmp(20256) := x"0000";
    tmp(20257) := x"0000";
    tmp(20258) := x"0020";
    tmp(20259) := x"0841";
    tmp(20260) := x"3986";
    tmp(20261) := x"628b";
    tmp(20262) := x"7aec";
    tmp(20263) := x"82cb";
    tmp(20264) := x"930b";
    tmp(20265) := x"8acb";
    tmp(20266) := x"92cb";
    tmp(20267) := x"bb4d";
    tmp(20268) := x"b2eb";
    tmp(20269) := x"d3ce";
    tmp(20270) := x"f532";
    tmp(20271) := x"a3ee";
    tmp(20272) := x"0841";
    tmp(20273) := x"0000";
    tmp(20274) := x"1040";
    tmp(20275) := x"8ae7";
    tmp(20276) := x"d48e";
    tmp(20277) := x"ab8c";
    tmp(20278) := x"938d";
    tmp(20279) := x"0000";
    tmp(20280) := x"20a1";
    tmp(20281) := x"f593";
    tmp(20282) := x"ab8e";
    tmp(20283) := x"938e";
    tmp(20284) := x"18a2";
    tmp(20285) := x"1061";
    tmp(20286) := x"1882";
    tmp(20287) := x"51a6";
    tmp(20288) := x"6a49";
    tmp(20289) := x"3124";
    tmp(20290) := x"1882";
    tmp(20291) := x"1061";
    tmp(20292) := x"0841";
    tmp(20293) := x"1041";
    tmp(20294) := x"20a2";
    tmp(20295) := x"5a06";
    tmp(20296) := x"3163";
    tmp(20297) := x"0040";
    tmp(20298) := x"08a0";
    tmp(20299) := x"08c0";
    tmp(20300) := x"08e0";
    tmp(20301) := x"0900";
    tmp(20302) := x"1140";
    tmp(20303) := x"1180";
    tmp(20304) := x"11a0";
    tmp(20305) := x"1a20";
    tmp(20306) := x"11e1";
    tmp(20307) := x"1a22";
    tmp(20308) := x"2b66";
    tmp(20309) := x"32c4";
    tmp(20310) := x"7447";
    tmp(20311) := x"9c69";
    tmp(20312) := x"ac8a";
    tmp(20313) := x"bccc";
    tmp(20314) := x"cd4d";
    tmp(20315) := x"ddaf";
    tmp(20316) := x"e630";
    tmp(20317) := x"e630";
    tmp(20318) := x"e610";
    tmp(20319) := x"e62f";
    tmp(20320) := x"d5ee";
    tmp(20321) := x"c58c";
    tmp(20322) := x"b50b";
    tmp(20323) := x"a48a";
    tmp(20324) := x"9c49";
    tmp(20325) := x"83a7";
    tmp(20326) := x"7b66";
    tmp(20327) := x"62e4";
    tmp(20328) := x"5283";
    tmp(20329) := x"4222";
    tmp(20330) := x"31c1";
    tmp(20331) := x"2961";
    tmp(20332) := x"2141";
    tmp(20333) := x"2981";
    tmp(20334) := x"31c2";
    tmp(20335) := x"39e3";
    tmp(20336) := x"4224";
    tmp(20337) := x"4a25";
    tmp(20338) := x"5246";
    tmp(20339) := x"5a67";
    tmp(20340) := x"6ae8";
    tmp(20341) := x"72e9";
    tmp(20342) := x"7b0a";
    tmp(20343) := x"834a";
    tmp(20344) := x"836a";
    tmp(20345) := x"7b4a";
    tmp(20346) := x"7b4a";
    tmp(20347) := x"836b";
    tmp(20348) := x"7b4a";
    tmp(20349) := x"7b6b";
    tmp(20350) := x"734b";
    tmp(20351) := x"736b";
    tmp(20352) := x"6b6a";
    tmp(20353) := x"6b2a";
    tmp(20354) := x"630a";
    tmp(20355) := x"632a";
    tmp(20356) := x"52a9";
    tmp(20357) := x"f800";
    tmp(20358) := x"f800";
    tmp(20359) := x"f800";
    tmp(20360) := x"f800";
    tmp(20361) := x"f800";
    tmp(20362) := x"f800";
    tmp(20363) := x"f800";
    tmp(20364) := x"f800";
    tmp(20365) := x"f800";
    tmp(20366) := x"f800";
    tmp(20367) := x"f800";
    tmp(20368) := x"f800";
    tmp(20369) := x"f800";
    tmp(20370) := x"f800";
    tmp(20371) := x"f800";
    tmp(20372) := x"f800";
    tmp(20373) := x"f800";
    tmp(20374) := x"f800";
    tmp(20375) := x"f800";
    tmp(20376) := x"f800";
    tmp(20377) := x"f800";
    tmp(20378) := x"f800";
    tmp(20379) := x"f800";
    tmp(20380) := x"f800";
    tmp(20381) := x"f800";
    tmp(20382) := x"f800";
    tmp(20383) := x"f800";
    tmp(20384) := x"f800";
    tmp(20385) := x"f800";
    tmp(20386) := x"f800";
    tmp(20387) := x"f800";
    tmp(20388) := x"f800";
    tmp(20389) := x"f800";
    tmp(20390) := x"f800";
    tmp(20391) := x"f800";
    tmp(20392) := x"f800";
    tmp(20393) := x"f800";
    tmp(20394) := x"f800";
    tmp(20395) := x"f800";
    tmp(20396) := x"f800";
    tmp(20397) := x"0840";
    tmp(20398) := x"0840";
    tmp(20399) := x"0840";
    tmp(20400) := x"1840";
    tmp(20401) := x"eb40";
    tmp(20402) := x"e300";
    tmp(20403) := x"e320";
    tmp(20404) := x"f340";
    tmp(20405) := x"f340";
    tmp(20406) := x"fb60";
    tmp(20407) := x"f340";
    tmp(20408) := x"f340";
    tmp(20409) := x"fb60";
    tmp(20410) := x"f360";
    tmp(20411) := x"f340";
    tmp(20412) := x"fba0";
    tmp(20413) := x"fb80";
    tmp(20414) := x"fba0";
    tmp(20415) := x"eb40";
    tmp(20416) := x"d300";
    tmp(20417) := x"c2e0";
    tmp(20418) := x"db20";
    tmp(20419) := x"d300";
    tmp(20420) := x"cae0";
    tmp(20421) := x"cae0";
    tmp(20422) := x"d300";
    tmp(20423) := x"db20";
    tmp(20424) := x"d300";
    tmp(20425) := x"d2e0";
    tmp(20426) := x"d300";
    tmp(20427) := x"d300";
    tmp(20428) := x"e340";
    tmp(20429) := x"f380";
    tmp(20430) := x"eb80";
    tmp(20431) := x"eb60";
    tmp(20432) := x"eba0";
    tmp(20433) := x"eb60";
    tmp(20434) := x"eb60";
    tmp(20435) := x"f380";
    tmp(20436) := x"f380";
    tmp(20437) := x"f360";
    tmp(20438) := x"eb40";
    tmp(20439) := x"eb40";
    tmp(20440) := x"f340";
    tmp(20441) := x"eb40";
    tmp(20442) := x"f360";
    tmp(20443) := x"fb80";
    tmp(20444) := x"fb60";
    tmp(20445) := x"fba0";
    tmp(20446) := x"fbc0";
    tmp(20447) := x"f360";
    tmp(20448) := x"cac0";
    tmp(20449) := x"c2c0";
    tmp(20450) := x"b260";
    tmp(20451) := x"ba60";
    tmp(20452) := x"c260";
    tmp(20453) := x"caa0";
    tmp(20454) := x"d2e0";
    tmp(20455) := x"e320";
    tmp(20456) := x"e340";
    tmp(20457) := x"d300";
    tmp(20458) := x"c2c0";
    tmp(20459) := x"baa0";
    tmp(20460) := x"b260";
    tmp(20461) := x"aa40";
    tmp(20462) := x"aa40";
    tmp(20463) := x"b260";
    tmp(20464) := x"b260";
    tmp(20465) := x"b260";
    tmp(20466) := x"aa40";
    tmp(20467) := x"aa40";
    tmp(20468) := x"b260";
    tmp(20469) := x"aa40";
    tmp(20470) := x"81c0";
    tmp(20471) := x"7180";
    tmp(20472) := x"6160";
    tmp(20473) := x"5140";
    tmp(20474) := x"3100";
    tmp(20475) := x"20a0";
    tmp(20476) := x"18a0";
    tmp(20477) := x"1080";
    tmp(20478) := x"0860";
    tmp(20479) := x"0860";
    tmp(20480) := x"0020";
    tmp(20481) := x"0000";
    tmp(20482) := x"0000";
    tmp(20483) := x"0020";
    tmp(20484) := x"0020";
    tmp(20485) := x"0020";
    tmp(20486) := x"0820";
    tmp(20487) := x"0820";
    tmp(20488) := x"0020";
    tmp(20489) := x"0000";
    tmp(20490) := x"0000";
    tmp(20491) := x"0000";
    tmp(20492) := x"0000";
    tmp(20493) := x"0000";
    tmp(20494) := x"0000";
    tmp(20495) := x"0000";
    tmp(20496) := x"0000";
    tmp(20497) := x"0000";
    tmp(20498) := x"0000";
    tmp(20499) := x"0000";
    tmp(20500) := x"0000";
    tmp(20501) := x"0000";
    tmp(20502) := x"0000";
    tmp(20503) := x"0020";
    tmp(20504) := x"0841";
    tmp(20505) := x"20c3";
    tmp(20506) := x"830c";
    tmp(20507) := x"7a8a";
    tmp(20508) := x"930c";
    tmp(20509) := x"72a9";
    tmp(20510) := x"20a2";
    tmp(20511) := x"0000";
    tmp(20512) := x"0000";
    tmp(20513) := x"1860";
    tmp(20514) := x"8ac2";
    tmp(20515) := x"69c2";
    tmp(20516) := x"28a0";
    tmp(20517) := x"a36a";
    tmp(20518) := x"0820";
    tmp(20519) := x"0000";
    tmp(20520) := x"8aea";
    tmp(20521) := x"bc10";
    tmp(20522) := x"9b6e";
    tmp(20523) := x"3145";
    tmp(20524) := x"0820";
    tmp(20525) := x"6aa9";
    tmp(20526) := x"5a28";
    tmp(20527) := x"3925";
    tmp(20528) := x"61e8";
    tmp(20529) := x"72ab";
    tmp(20530) := x"5208";
    tmp(20531) := x"41a6";
    tmp(20532) := x"3985";
    tmp(20533) := x"3964";
    tmp(20534) := x"20e2";
    tmp(20535) := x"1081";
    tmp(20536) := x"0840";
    tmp(20537) := x"0880";
    tmp(20538) := x"08c0";
    tmp(20539) := x"08c0";
    tmp(20540) := x"08c0";
    tmp(20541) := x"1120";
    tmp(20542) := x"1160";
    tmp(20543) := x"19c0";
    tmp(20544) := x"11c0";
    tmp(20545) := x"1a21";
    tmp(20546) := x"1aa2";
    tmp(20547) := x"1a42";
    tmp(20548) := x"3c06";
    tmp(20549) := x"6c48";
    tmp(20550) := x"73a7";
    tmp(20551) := x"93e8";
    tmp(20552) := x"a44a";
    tmp(20553) := x"bccb";
    tmp(20554) := x"cd6d";
    tmp(20555) := x"ddaf";
    tmp(20556) := x"ddf0";
    tmp(20557) := x"e631";
    tmp(20558) := x"e610";
    tmp(20559) := x"e650";
    tmp(20560) := x"ee6f";
    tmp(20561) := x"de0e";
    tmp(20562) := x"ddee";
    tmp(20563) := x"c56d";
    tmp(20564) := x"b4cb";
    tmp(20565) := x"a4aa";
    tmp(20566) := x"9428";
    tmp(20567) := x"7b86";
    tmp(20568) := x"6b25";
    tmp(20569) := x"5ac4";
    tmp(20570) := x"4a42";
    tmp(20571) := x"39e2";
    tmp(20572) := x"2981";
    tmp(20573) := x"2961";
    tmp(20574) := x"29a2";
    tmp(20575) := x"39e3";
    tmp(20576) := x"3a04";
    tmp(20577) := x"4a45";
    tmp(20578) := x"5266";
    tmp(20579) := x"5a87";
    tmp(20580) := x"6ac8";
    tmp(20581) := x"7309";
    tmp(20582) := x"7b2a";
    tmp(20583) := x"7b4a";
    tmp(20584) := x"834b";
    tmp(20585) := x"8b6c";
    tmp(20586) := x"8b6c";
    tmp(20587) := x"8b6b";
    tmp(20588) := x"8b8c";
    tmp(20589) := x"836c";
    tmp(20590) := x"7b6b";
    tmp(20591) := x"838c";
    tmp(20592) := x"7bac";
    tmp(20593) := x"6b4b";
    tmp(20594) := x"6b2b";
    tmp(20595) := x"632b";
    tmp(20596) := x"5aea";
    tmp(20597) := x"f800";
    tmp(20598) := x"f800";
    tmp(20599) := x"f800";
    tmp(20600) := x"f800";
    tmp(20601) := x"f800";
    tmp(20602) := x"f800";
    tmp(20603) := x"f800";
    tmp(20604) := x"f800";
    tmp(20605) := x"f800";
    tmp(20606) := x"f800";
    tmp(20607) := x"f800";
    tmp(20608) := x"f800";
    tmp(20609) := x"f800";
    tmp(20610) := x"f800";
    tmp(20611) := x"f800";
    tmp(20612) := x"f800";
    tmp(20613) := x"f800";
    tmp(20614) := x"f800";
    tmp(20615) := x"f800";
    tmp(20616) := x"f800";
    tmp(20617) := x"f800";
    tmp(20618) := x"f800";
    tmp(20619) := x"f800";
    tmp(20620) := x"f800";
    tmp(20621) := x"f800";
    tmp(20622) := x"f800";
    tmp(20623) := x"f800";
    tmp(20624) := x"f800";
    tmp(20625) := x"f800";
    tmp(20626) := x"f800";
    tmp(20627) := x"f800";
    tmp(20628) := x"f800";
    tmp(20629) := x"f800";
    tmp(20630) := x"f800";
    tmp(20631) := x"f800";
    tmp(20632) := x"f800";
    tmp(20633) := x"f800";
    tmp(20634) := x"f800";
    tmp(20635) := x"f800";
    tmp(20636) := x"f800";
    tmp(20637) := x"0840";
    tmp(20638) := x"0840";
    tmp(20639) := x"0840";
    tmp(20640) := x"1840";
    tmp(20641) := x"eb40";
    tmp(20642) := x"db20";
    tmp(20643) := x"e340";
    tmp(20644) := x"eb20";
    tmp(20645) := x"eb20";
    tmp(20646) := x"fb40";
    tmp(20647) := x"f340";
    tmp(20648) := x"fb80";
    tmp(20649) := x"fb60";
    tmp(20650) := x"fb80";
    tmp(20651) := x"f360";
    tmp(20652) := x"fba0";
    tmp(20653) := x"fba0";
    tmp(20654) := x"fba0";
    tmp(20655) := x"eb80";
    tmp(20656) := x"eb60";
    tmp(20657) := x"db40";
    tmp(20658) := x"c2e0";
    tmp(20659) := x"ba80";
    tmp(20660) := x"cac0";
    tmp(20661) := x"db00";
    tmp(20662) := x"db20";
    tmp(20663) := x"db20";
    tmp(20664) := x"d320";
    tmp(20665) := x"d300";
    tmp(20666) := x"d2e0";
    tmp(20667) := x"db20";
    tmp(20668) := x"db00";
    tmp(20669) := x"fba0";
    tmp(20670) := x"e340";
    tmp(20671) := x"f380";
    tmp(20672) := x"fbc0";
    tmp(20673) := x"f360";
    tmp(20674) := x"eb60";
    tmp(20675) := x"fb80";
    tmp(20676) := x"fba0";
    tmp(20677) := x"f380";
    tmp(20678) := x"f340";
    tmp(20679) := x"f340";
    tmp(20680) := x"eb40";
    tmp(20681) := x"f360";
    tmp(20682) := x"fb80";
    tmp(20683) := x"f360";
    tmp(20684) := x"fb60";
    tmp(20685) := x"fb80";
    tmp(20686) := x"fba0";
    tmp(20687) := x"fb80";
    tmp(20688) := x"eb20";
    tmp(20689) := x"c280";
    tmp(20690) := x"ba60";
    tmp(20691) := x"ba40";
    tmp(20692) := x"c260";
    tmp(20693) := x"caa0";
    tmp(20694) := x"dae0";
    tmp(20695) := x"d2e0";
    tmp(20696) := x"db20";
    tmp(20697) := x"cb00";
    tmp(20698) := x"c2e0";
    tmp(20699) := x"c2e0";
    tmp(20700) := x"aa80";
    tmp(20701) := x"ba80";
    tmp(20702) := x"b280";
    tmp(20703) := x"ba80";
    tmp(20704) := x"ba80";
    tmp(20705) := x"ba80";
    tmp(20706) := x"ba80";
    tmp(20707) := x"b260";
    tmp(20708) := x"aa40";
    tmp(20709) := x"aa40";
    tmp(20710) := x"b280";
    tmp(20711) := x"b280";
    tmp(20712) := x"9a20";
    tmp(20713) := x"89e0";
    tmp(20714) := x"6180";
    tmp(20715) := x"4120";
    tmp(20716) := x"28c0";
    tmp(20717) := x"1080";
    tmp(20718) := x"0860";
    tmp(20719) := x"0840";
    tmp(20720) := x"0820";
    tmp(20721) := x"0020";
    tmp(20722) := x"0000";
    tmp(20723) := x"0020";
    tmp(20724) := x"0020";
    tmp(20725) := x"0840";
    tmp(20726) := x"0820";
    tmp(20727) := x"0820";
    tmp(20728) := x"0020";
    tmp(20729) := x"0000";
    tmp(20730) := x"0000";
    tmp(20731) := x"0000";
    tmp(20732) := x"0000";
    tmp(20733) := x"0000";
    tmp(20734) := x"0000";
    tmp(20735) := x"0000";
    tmp(20736) := x"0000";
    tmp(20737) := x"0000";
    tmp(20738) := x"0000";
    tmp(20739) := x"0000";
    tmp(20740) := x"0000";
    tmp(20741) := x"0000";
    tmp(20742) := x"0000";
    tmp(20743) := x"0020";
    tmp(20744) := x"0000";
    tmp(20745) := x"0000";
    tmp(20746) := x"0000";
    tmp(20747) := x"0821";
    tmp(20748) := x"0841";
    tmp(20749) := x"0000";
    tmp(20750) := x"0000";
    tmp(20751) := x"0820";
    tmp(20752) := x"28c0";
    tmp(20753) := x"69c0";
    tmp(20754) := x"38e0";
    tmp(20755) := x"2080";
    tmp(20756) := x"59a1";
    tmp(20757) := x"3102";
    tmp(20758) := x"0000";
    tmp(20759) := x"3943";
    tmp(20760) := x"cc91";
    tmp(20761) := x"8b2c";
    tmp(20762) := x"3965";
    tmp(20763) := x"0000";
    tmp(20764) := x"1881";
    tmp(20765) := x"dd33";
    tmp(20766) := x"932d";
    tmp(20767) := x"7a8a";
    tmp(20768) := x"728a";
    tmp(20769) := x"51c7";
    tmp(20770) := x"41c6";
    tmp(20771) := x"2103";
    tmp(20772) := x"1081";
    tmp(20773) := x"0840";
    tmp(20774) := x"0040";
    tmp(20775) := x"0860";
    tmp(20776) := x"0880";
    tmp(20777) := x"08a0";
    tmp(20778) := x"08c0";
    tmp(20779) := x"08c0";
    tmp(20780) := x"1120";
    tmp(20781) := x"1140";
    tmp(20782) := x"1180";
    tmp(20783) := x"19e0";
    tmp(20784) := x"1a21";
    tmp(20785) := x"1a02";
    tmp(20786) := x"11e1";
    tmp(20787) := x"3383";
    tmp(20788) := x"4c06";
    tmp(20789) := x"52e5";
    tmp(20790) := x"6b46";
    tmp(20791) := x"83a7";
    tmp(20792) := x"9409";
    tmp(20793) := x"ac8a";
    tmp(20794) := x"bcec";
    tmp(20795) := x"cd6d";
    tmp(20796) := x"ddef";
    tmp(20797) := x"ee30";
    tmp(20798) := x"f691";
    tmp(20799) := x"f6b1";
    tmp(20800) := x"ee50";
    tmp(20801) := x"f691";
    tmp(20802) := x"ee70";
    tmp(20803) := x"e66f";
    tmp(20804) := x"d5ee";
    tmp(20805) := x"bd6c";
    tmp(20806) := x"acca";
    tmp(20807) := x"9c69";
    tmp(20808) := x"83c7";
    tmp(20809) := x"7346";
    tmp(20810) := x"5ac4";
    tmp(20811) := x"5263";
    tmp(20812) := x"4202";
    tmp(20813) := x"31c1";
    tmp(20814) := x"31a2";
    tmp(20815) := x"31a2";
    tmp(20816) := x"4224";
    tmp(20817) := x"4a45";
    tmp(20818) := x"4a65";
    tmp(20819) := x"5a86";
    tmp(20820) := x"62a7";
    tmp(20821) := x"7309";
    tmp(20822) := x"7b4a";
    tmp(20823) := x"834b";
    tmp(20824) := x"8b6c";
    tmp(20825) := x"93ad";
    tmp(20826) := x"93ad";
    tmp(20827) := x"93ad";
    tmp(20828) := x"8bad";
    tmp(20829) := x"93cd";
    tmp(20830) := x"8bad";
    tmp(20831) := x"8bcd";
    tmp(20832) := x"8bcd";
    tmp(20833) := x"7bad";
    tmp(20834) := x"7b6d";
    tmp(20835) := x"6b4c";
    tmp(20836) := x"630b";
    tmp(20837) := x"f800";
    tmp(20838) := x"f800";
    tmp(20839) := x"f800";
    tmp(20840) := x"f800";
    tmp(20841) := x"f800";
    tmp(20842) := x"f800";
    tmp(20843) := x"f800";
    tmp(20844) := x"f800";
    tmp(20845) := x"f800";
    tmp(20846) := x"f800";
    tmp(20847) := x"f800";
    tmp(20848) := x"f800";
    tmp(20849) := x"f800";
    tmp(20850) := x"f800";
    tmp(20851) := x"f800";
    tmp(20852) := x"f800";
    tmp(20853) := x"f800";
    tmp(20854) := x"f800";
    tmp(20855) := x"f800";
    tmp(20856) := x"f800";
    tmp(20857) := x"f800";
    tmp(20858) := x"f800";
    tmp(20859) := x"f800";
    tmp(20860) := x"f800";
    tmp(20861) := x"f800";
    tmp(20862) := x"f800";
    tmp(20863) := x"f800";
    tmp(20864) := x"f800";
    tmp(20865) := x"f800";
    tmp(20866) := x"f800";
    tmp(20867) := x"f800";
    tmp(20868) := x"f800";
    tmp(20869) := x"f800";
    tmp(20870) := x"f800";
    tmp(20871) := x"f800";
    tmp(20872) := x"f800";
    tmp(20873) := x"f800";
    tmp(20874) := x"f800";
    tmp(20875) := x"f800";
    tmp(20876) := x"f800";
    tmp(20877) := x"0840";
    tmp(20878) := x"0840";
    tmp(20879) := x"0840";
    tmp(20880) := x"1040";
    tmp(20881) := x"f360";
    tmp(20882) := x"e340";
    tmp(20883) := x"e320";
    tmp(20884) := x"eb20";
    tmp(20885) := x"f340";
    tmp(20886) := x"fb60";
    tmp(20887) := x"fb60";
    tmp(20888) := x"f360";
    tmp(20889) := x"f380";
    tmp(20890) := x"f360";
    tmp(20891) := x"fb80";
    tmp(20892) := x"f380";
    tmp(20893) := x"fba0";
    tmp(20894) := x"fb80";
    tmp(20895) := x"f380";
    tmp(20896) := x"eb80";
    tmp(20897) := x"d320";
    tmp(20898) := x"cb00";
    tmp(20899) := x"cac0";
    tmp(20900) := x"db20";
    tmp(20901) := x"d2e0";
    tmp(20902) := x"d2e0";
    tmp(20903) := x"cae0";
    tmp(20904) := x"cac0";
    tmp(20905) := x"d300";
    tmp(20906) := x"d2e0";
    tmp(20907) := x"db20";
    tmp(20908) := x"db40";
    tmp(20909) := x"e340";
    tmp(20910) := x"e340";
    tmp(20911) := x"eb60";
    tmp(20912) := x"fba0";
    tmp(20913) := x"eb60";
    tmp(20914) := x"f340";
    tmp(20915) := x"f340";
    tmp(20916) := x"f340";
    tmp(20917) := x"f340";
    tmp(20918) := x"fb40";
    tmp(20919) := x"f340";
    tmp(20920) := x"fb60";
    tmp(20921) := x"eb40";
    tmp(20922) := x"fb60";
    tmp(20923) := x"fb80";
    tmp(20924) := x"fb60";
    tmp(20925) := x"fb40";
    tmp(20926) := x"eb40";
    tmp(20927) := x"f360";
    tmp(20928) := x"f360";
    tmp(20929) := x"dae0";
    tmp(20930) := x"d2a0";
    tmp(20931) := x"caa0";
    tmp(20932) := x"caa0";
    tmp(20933) := x"caa0";
    tmp(20934) := x"dae0";
    tmp(20935) := x"e320";
    tmp(20936) := x"db20";
    tmp(20937) := x"d320";
    tmp(20938) := x"d320";
    tmp(20939) := x"cae0";
    tmp(20940) := x"baa0";
    tmp(20941) := x"c2c0";
    tmp(20942) := x"c2c0";
    tmp(20943) := x"baa0";
    tmp(20944) := x"c2a0";
    tmp(20945) := x"baa0";
    tmp(20946) := x"b280";
    tmp(20947) := x"b260";
    tmp(20948) := x"aa40";
    tmp(20949) := x"b240";
    tmp(20950) := x"ba80";
    tmp(20951) := x"ba80";
    tmp(20952) := x"b260";
    tmp(20953) := x"9200";
    tmp(20954) := x"81e0";
    tmp(20955) := x"5960";
    tmp(20956) := x"38e0";
    tmp(20957) := x"18a0";
    tmp(20958) := x"0860";
    tmp(20959) := x"0860";
    tmp(20960) := x"0840";
    tmp(20961) := x"0020";
    tmp(20962) := x"0020";
    tmp(20963) := x"0020";
    tmp(20964) := x"0020";
    tmp(20965) := x"0840";
    tmp(20966) := x"0840";
    tmp(20967) := x"0840";
    tmp(20968) := x"0020";
    tmp(20969) := x"0020";
    tmp(20970) := x"0000";
    tmp(20971) := x"0000";
    tmp(20972) := x"0000";
    tmp(20973) := x"0000";
    tmp(20974) := x"0000";
    tmp(20975) := x"0000";
    tmp(20976) := x"0000";
    tmp(20977) := x"0000";
    tmp(20978) := x"0000";
    tmp(20979) := x"0000";
    tmp(20980) := x"0000";
    tmp(20981) := x"0820";
    tmp(20982) := x"0820";
    tmp(20983) := x"0000";
    tmp(20984) := x"0000";
    tmp(20985) := x"0000";
    tmp(20986) := x"0000";
    tmp(20987) := x"0000";
    tmp(20988) := x"0000";
    tmp(20989) := x"0020";
    tmp(20990) := x"0840";
    tmp(20991) := x"30e0";
    tmp(20992) := x"5160";
    tmp(20993) := x"28c0";
    tmp(20994) := x"20a0";
    tmp(20995) := x"4120";
    tmp(20996) := x"59e2";
    tmp(20997) := x"0020";
    tmp(20998) := x"0840";
    tmp(20999) := x"bc8e";
    tmp(21000) := x"6248";
    tmp(21001) := x"1882";
    tmp(21002) := x"0000";
    tmp(21003) := x"0820";
    tmp(21004) := x"8b4b";
    tmp(21005) := x"bc10";
    tmp(21006) := x"bc52";
    tmp(21007) := x"936d";
    tmp(21008) := x"6ac9";
    tmp(21009) := x"39c4";
    tmp(21010) := x"10a1";
    tmp(21011) := x"0880";
    tmp(21012) := x"0860";
    tmp(21013) := x"08a0";
    tmp(21014) := x"08a0";
    tmp(21015) := x"08a0";
    tmp(21016) := x"08c0";
    tmp(21017) := x"08c0";
    tmp(21018) := x"08e0";
    tmp(21019) := x"1140";
    tmp(21020) := x"1140";
    tmp(21021) := x"11a0";
    tmp(21022) := x"1a01";
    tmp(21023) := x"2241";
    tmp(21024) := x"1a02";
    tmp(21025) := x"1a01";
    tmp(21026) := x"1a42";
    tmp(21027) := x"43e5";
    tmp(21028) := x"3a43";
    tmp(21029) := x"4a63";
    tmp(21030) := x"62e5";
    tmp(21031) := x"7366";
    tmp(21032) := x"8bc7";
    tmp(21033) := x"a46a";
    tmp(21034) := x"b4ab";
    tmp(21035) := x"c54d";
    tmp(21036) := x"ddef";
    tmp(21037) := x"e60f";
    tmp(21038) := x"f670";
    tmp(21039) := x"fed2";
    tmp(21040) := x"fef2";
    tmp(21041) := x"ff13";
    tmp(21042) := x"fed2";
    tmp(21043) := x"f6b1";
    tmp(21044) := x"f691";
    tmp(21045) := x"de2f";
    tmp(21046) := x"cdad";
    tmp(21047) := x"b50b";
    tmp(21048) := x"a469";
    tmp(21049) := x"8be8";
    tmp(21050) := x"7b46";
    tmp(21051) := x"62e5";
    tmp(21052) := x"5283";
    tmp(21053) := x"4202";
    tmp(21054) := x"39c2";
    tmp(21055) := x"31a2";
    tmp(21056) := x"3a03";
    tmp(21057) := x"4224";
    tmp(21058) := x"5265";
    tmp(21059) := x"5a86";
    tmp(21060) := x"62c8";
    tmp(21061) := x"6ae9";
    tmp(21062) := x"7b2a";
    tmp(21063) := x"8b6c";
    tmp(21064) := x"8b8d";
    tmp(21065) := x"93ad";
    tmp(21066) := x"9bce";
    tmp(21067) := x"9bee";
    tmp(21068) := x"9bef";
    tmp(21069) := x"9c0f";
    tmp(21070) := x"940f";
    tmp(21071) := x"942e";
    tmp(21072) := x"8bee";
    tmp(21073) := x"8bee";
    tmp(21074) := x"83ce";
    tmp(21075) := x"736d";
    tmp(21076) := x"6b4c";
    tmp(21077) := x"f800";
    tmp(21078) := x"f800";
    tmp(21079) := x"f800";
    tmp(21080) := x"f800";
    tmp(21081) := x"f800";
    tmp(21082) := x"f800";
    tmp(21083) := x"f800";
    tmp(21084) := x"f800";
    tmp(21085) := x"f800";
    tmp(21086) := x"f800";
    tmp(21087) := x"f800";
    tmp(21088) := x"f800";
    tmp(21089) := x"f800";
    tmp(21090) := x"f800";
    tmp(21091) := x"f800";
    tmp(21092) := x"f800";
    tmp(21093) := x"f800";
    tmp(21094) := x"f800";
    tmp(21095) := x"f800";
    tmp(21096) := x"f800";
    tmp(21097) := x"f800";
    tmp(21098) := x"f800";
    tmp(21099) := x"f800";
    tmp(21100) := x"f800";
    tmp(21101) := x"f800";
    tmp(21102) := x"f800";
    tmp(21103) := x"f800";
    tmp(21104) := x"f800";
    tmp(21105) := x"f800";
    tmp(21106) := x"f800";
    tmp(21107) := x"f800";
    tmp(21108) := x"f800";
    tmp(21109) := x"f800";
    tmp(21110) := x"f800";
    tmp(21111) := x"f800";
    tmp(21112) := x"f800";
    tmp(21113) := x"f800";
    tmp(21114) := x"f800";
    tmp(21115) := x"f800";
    tmp(21116) := x"f800";
    tmp(21117) := x"0840";
    tmp(21118) := x"0840";
    tmp(21119) := x"0840";
    tmp(21120) := x"1040";
    tmp(21121) := x"eb60";
    tmp(21122) := x"db20";
    tmp(21123) := x"eb40";
    tmp(21124) := x"f340";
    tmp(21125) := x"f360";
    tmp(21126) := x"fb60";
    tmp(21127) := x"fb60";
    tmp(21128) := x"fb80";
    tmp(21129) := x"f360";
    tmp(21130) := x"f380";
    tmp(21131) := x"fba0";
    tmp(21132) := x"fba0";
    tmp(21133) := x"fba0";
    tmp(21134) := x"fb80";
    tmp(21135) := x"fba0";
    tmp(21136) := x"f380";
    tmp(21137) := x"db20";
    tmp(21138) := x"d300";
    tmp(21139) := x"d2e0";
    tmp(21140) := x"d2e0";
    tmp(21141) := x"d2c0";
    tmp(21142) := x"d2c0";
    tmp(21143) := x"d2c0";
    tmp(21144) := x"cac0";
    tmp(21145) := x"cac0";
    tmp(21146) := x"d2c0";
    tmp(21147) := x"db00";
    tmp(21148) := x"db00";
    tmp(21149) := x"f360";
    tmp(21150) := x"eb40";
    tmp(21151) := x"e340";
    tmp(21152) := x"eb60";
    tmp(21153) := x"f340";
    tmp(21154) := x"eb20";
    tmp(21155) := x"f340";
    tmp(21156) := x"fb60";
    tmp(21157) := x"f360";
    tmp(21158) := x"f340";
    tmp(21159) := x"f360";
    tmp(21160) := x"fb60";
    tmp(21161) := x"fb60";
    tmp(21162) := x"eb40";
    tmp(21163) := x"fb40";
    tmp(21164) := x"fb40";
    tmp(21165) := x"eb20";
    tmp(21166) := x"fba0";
    tmp(21167) := x"fba0";
    tmp(21168) := x"f380";
    tmp(21169) := x"eb40";
    tmp(21170) := x"dae0";
    tmp(21171) := x"d2c0";
    tmp(21172) := x"d2a0";
    tmp(21173) := x"dac0";
    tmp(21174) := x"dac0";
    tmp(21175) := x"dae0";
    tmp(21176) := x"db20";
    tmp(21177) := x"d300";
    tmp(21178) := x"cae0";
    tmp(21179) := x"baa0";
    tmp(21180) := x"c2c0";
    tmp(21181) := x"baa0";
    tmp(21182) := x"c2c0";
    tmp(21183) := x"c2c0";
    tmp(21184) := x"c2c0";
    tmp(21185) := x"c2a0";
    tmp(21186) := x"ba80";
    tmp(21187) := x"ba80";
    tmp(21188) := x"c2a0";
    tmp(21189) := x"ba60";
    tmp(21190) := x"b240";
    tmp(21191) := x"ba40";
    tmp(21192) := x"ba60";
    tmp(21193) := x"b260";
    tmp(21194) := x"9a20";
    tmp(21195) := x"81e0";
    tmp(21196) := x"5960";
    tmp(21197) := x"30e0";
    tmp(21198) := x"1080";
    tmp(21199) := x"0840";
    tmp(21200) := x"0020";
    tmp(21201) := x"0840";
    tmp(21202) := x"0020";
    tmp(21203) := x"0020";
    tmp(21204) := x"0020";
    tmp(21205) := x"0840";
    tmp(21206) := x"0840";
    tmp(21207) := x"0840";
    tmp(21208) := x"0020";
    tmp(21209) := x"0020";
    tmp(21210) := x"0020";
    tmp(21211) := x"0000";
    tmp(21212) := x"0000";
    tmp(21213) := x"0000";
    tmp(21214) := x"0000";
    tmp(21215) := x"0000";
    tmp(21216) := x"0000";
    tmp(21217) := x"0020";
    tmp(21218) := x"0020";
    tmp(21219) := x"0820";
    tmp(21220) := x"0820";
    tmp(21221) := x"0820";
    tmp(21222) := x"0020";
    tmp(21223) := x"0000";
    tmp(21224) := x"0000";
    tmp(21225) := x"0000";
    tmp(21226) := x"0000";
    tmp(21227) := x"0000";
    tmp(21228) := x"0820";
    tmp(21229) := x"1060";
    tmp(21230) := x"3900";
    tmp(21231) := x"5140";
    tmp(21232) := x"30e0";
    tmp(21233) := x"28c0";
    tmp(21234) := x"4940";
    tmp(21235) := x"69c0";
    tmp(21236) := x"1060";
    tmp(21237) := x"0820";
    tmp(21238) := x"20a1";
    tmp(21239) := x"3143";
    tmp(21240) := x"0000";
    tmp(21241) := x"0000";
    tmp(21242) := x"0840";
    tmp(21243) := x"49c5";
    tmp(21244) := x"b40f";
    tmp(21245) := x"9b6d";
    tmp(21246) := x"834b";
    tmp(21247) := x"4205";
    tmp(21248) := x"18e1";
    tmp(21249) := x"0860";
    tmp(21250) := x"0860";
    tmp(21251) := x"0880";
    tmp(21252) := x"08a0";
    tmp(21253) := x"08c0";
    tmp(21254) := x"08a0";
    tmp(21255) := x"08c0";
    tmp(21256) := x"08c0";
    tmp(21257) := x"0900";
    tmp(21258) := x"1140";
    tmp(21259) := x"1140";
    tmp(21260) := x"11c1";
    tmp(21261) := x"19e1";
    tmp(21262) := x"19e1";
    tmp(21263) := x"1a41";
    tmp(21264) := x"1a42";
    tmp(21265) := x"1a62";
    tmp(21266) := x"3344";
    tmp(21267) := x"29e2";
    tmp(21268) := x"31c2";
    tmp(21269) := x"4223";
    tmp(21270) := x"5263";
    tmp(21271) := x"6305";
    tmp(21272) := x"83a7";
    tmp(21273) := x"9c29";
    tmp(21274) := x"b4aa";
    tmp(21275) := x"bcec";
    tmp(21276) := x"cd6d";
    tmp(21277) := x"e5ee";
    tmp(21278) := x"f650";
    tmp(21279) := x"fed2";
    tmp(21280) := x"fef2";
    tmp(21281) := x"ff33";
    tmp(21282) := x"ff53";
    tmp(21283) := x"ff33";
    tmp(21284) := x"ff74";
    tmp(21285) := x"f6d2";
    tmp(21286) := x"ee90";
    tmp(21287) := x"ddee";
    tmp(21288) := x"c52c";
    tmp(21289) := x"b4ca";
    tmp(21290) := x"93e8";
    tmp(21291) := x"7b66";
    tmp(21292) := x"62e5";
    tmp(21293) := x"5aa4";
    tmp(21294) := x"4a43";
    tmp(21295) := x"39e2";
    tmp(21296) := x"39c2";
    tmp(21297) := x"3a03";
    tmp(21298) := x"4a65";
    tmp(21299) := x"5286";
    tmp(21300) := x"62c8";
    tmp(21301) := x"6b09";
    tmp(21302) := x"7b2a";
    tmp(21303) := x"7b4b";
    tmp(21304) := x"93ad";
    tmp(21305) := x"93ce";
    tmp(21306) := x"a3ef";
    tmp(21307) := x"a430";
    tmp(21308) := x"a410";
    tmp(21309) := x"a410";
    tmp(21310) := x"a451";
    tmp(21311) := x"9c71";
    tmp(21312) := x"9450";
    tmp(21313) := x"942f";
    tmp(21314) := x"8bcf";
    tmp(21315) := x"7b6e";
    tmp(21316) := x"732c";
    tmp(21317) := x"f800";
    tmp(21318) := x"f800";
    tmp(21319) := x"f800";
    tmp(21320) := x"f800";
    tmp(21321) := x"f800";
    tmp(21322) := x"f800";
    tmp(21323) := x"f800";
    tmp(21324) := x"f800";
    tmp(21325) := x"f800";
    tmp(21326) := x"f800";
    tmp(21327) := x"f800";
    tmp(21328) := x"f800";
    tmp(21329) := x"f800";
    tmp(21330) := x"f800";
    tmp(21331) := x"f800";
    tmp(21332) := x"f800";
    tmp(21333) := x"f800";
    tmp(21334) := x"f800";
    tmp(21335) := x"f800";
    tmp(21336) := x"f800";
    tmp(21337) := x"f800";
    tmp(21338) := x"f800";
    tmp(21339) := x"f800";
    tmp(21340) := x"f800";
    tmp(21341) := x"f800";
    tmp(21342) := x"f800";
    tmp(21343) := x"f800";
    tmp(21344) := x"f800";
    tmp(21345) := x"f800";
    tmp(21346) := x"f800";
    tmp(21347) := x"f800";
    tmp(21348) := x"f800";
    tmp(21349) := x"f800";
    tmp(21350) := x"f800";
    tmp(21351) := x"f800";
    tmp(21352) := x"f800";
    tmp(21353) := x"f800";
    tmp(21354) := x"f800";
    tmp(21355) := x"f800";
    tmp(21356) := x"f800";
    tmp(21357) := x"0840";
    tmp(21358) := x"0840";
    tmp(21359) := x"0840";
    tmp(21360) := x"1860";
    tmp(21361) := x"f340";
    tmp(21362) := x"e300";
    tmp(21363) := x"eb40";
    tmp(21364) := x"fb40";
    tmp(21365) := x"fb40";
    tmp(21366) := x"f340";
    tmp(21367) := x"fb40";
    tmp(21368) := x"fb60";
    tmp(21369) := x"f360";
    tmp(21370) := x"f360";
    tmp(21371) := x"fb80";
    tmp(21372) := x"fb80";
    tmp(21373) := x"fba0";
    tmp(21374) := x"fbc0";
    tmp(21375) := x"fbc0";
    tmp(21376) := x"fba0";
    tmp(21377) := x"eb40";
    tmp(21378) := x"db00";
    tmp(21379) := x"dae0";
    tmp(21380) := x"d2c0";
    tmp(21381) := x"dac0";
    tmp(21382) := x"e2e0";
    tmp(21383) := x"d2a0";
    tmp(21384) := x"caa0";
    tmp(21385) := x"cac0";
    tmp(21386) := x"d2c0";
    tmp(21387) := x"d2e0";
    tmp(21388) := x"dae0";
    tmp(21389) := x"e320";
    tmp(21390) := x"eb40";
    tmp(21391) := x"eb40";
    tmp(21392) := x"eb40";
    tmp(21393) := x"eb20";
    tmp(21394) := x"eb20";
    tmp(21395) := x"eb20";
    tmp(21396) := x"fb40";
    tmp(21397) := x"f360";
    tmp(21398) := x"f360";
    tmp(21399) := x"fb60";
    tmp(21400) := x"fb60";
    tmp(21401) := x"fb60";
    tmp(21402) := x"f340";
    tmp(21403) := x"f340";
    tmp(21404) := x"eb00";
    tmp(21405) := x"f340";
    tmp(21406) := x"fba0";
    tmp(21407) := x"fba0";
    tmp(21408) := x"fba0";
    tmp(21409) := x"f360";
    tmp(21410) := x"eb20";
    tmp(21411) := x"dae0";
    tmp(21412) := x"d2c0";
    tmp(21413) := x"dac0";
    tmp(21414) := x"dae0";
    tmp(21415) := x"e300";
    tmp(21416) := x"e320";
    tmp(21417) := x"e320";
    tmp(21418) := x"db00";
    tmp(21419) := x"c2a0";
    tmp(21420) := x"c2a0";
    tmp(21421) := x"c2a0";
    tmp(21422) := x"cb00";
    tmp(21423) := x"d300";
    tmp(21424) := x"cae0";
    tmp(21425) := x"cac0";
    tmp(21426) := x"cac0";
    tmp(21427) := x"cac0";
    tmp(21428) := x"cac0";
    tmp(21429) := x"ba60";
    tmp(21430) := x"b220";
    tmp(21431) := x"b240";
    tmp(21432) := x"ba40";
    tmp(21433) := x"c280";
    tmp(21434) := x"c280";
    tmp(21435) := x"aa40";
    tmp(21436) := x"8a00";
    tmp(21437) := x"5960";
    tmp(21438) := x"20a0";
    tmp(21439) := x"0840";
    tmp(21440) := x"0020";
    tmp(21441) := x"0020";
    tmp(21442) := x"0020";
    tmp(21443) := x"0040";
    tmp(21444) := x"0040";
    tmp(21445) := x"0840";
    tmp(21446) := x"0840";
    tmp(21447) := x"0840";
    tmp(21448) := x"0840";
    tmp(21449) := x"0020";
    tmp(21450) := x"0020";
    tmp(21451) := x"0000";
    tmp(21452) := x"0000";
    tmp(21453) := x"0000";
    tmp(21454) := x"0000";
    tmp(21455) := x"0000";
    tmp(21456) := x"0020";
    tmp(21457) := x"0840";
    tmp(21458) := x"1040";
    tmp(21459) := x"1040";
    tmp(21460) := x"1040";
    tmp(21461) := x"1040";
    tmp(21462) := x"1040";
    tmp(21463) := x"1040";
    tmp(21464) := x"0820";
    tmp(21465) := x"0000";
    tmp(21466) := x"0820";
    tmp(21467) := x"1040";
    tmp(21468) := x"28a0";
    tmp(21469) := x"5140";
    tmp(21470) := x"6960";
    tmp(21471) := x"4920";
    tmp(21472) := x"3900";
    tmp(21473) := x"5160";
    tmp(21474) := x"69a0";
    tmp(21475) := x"4940";
    tmp(21476) := x"0840";
    tmp(21477) := x"1080";
    tmp(21478) := x"3140";
    tmp(21479) := x"0000";
    tmp(21480) := x"0020";
    tmp(21481) := x"18a2";
    tmp(21482) := x"6a87";
    tmp(21483) := x"7b0a";
    tmp(21484) := x"5246";
    tmp(21485) := x"2963";
    tmp(21486) := x"10c1";
    tmp(21487) := x"0840";
    tmp(21488) := x"0060";
    tmp(21489) := x"0880";
    tmp(21490) := x"08a0";
    tmp(21491) := x"0880";
    tmp(21492) := x"0880";
    tmp(21493) := x"08c0";
    tmp(21494) := x"08c0";
    tmp(21495) := x"08c0";
    tmp(21496) := x"08e0";
    tmp(21497) := x"1140";
    tmp(21498) := x"0920";
    tmp(21499) := x"1181";
    tmp(21500) := x"1a02";
    tmp(21501) := x"11a1";
    tmp(21502) := x"1a21";
    tmp(21503) := x"22c3";
    tmp(21504) := x"2283";
    tmp(21505) := x"2ac3";
    tmp(21506) := x"21e2";
    tmp(21507) := x"2181";
    tmp(21508) := x"2981";
    tmp(21509) := x"31e2";
    tmp(21510) := x"4243";
    tmp(21511) := x"5ac4";
    tmp(21512) := x"7345";
    tmp(21513) := x"8bc8";
    tmp(21514) := x"a449";
    tmp(21515) := x"bceb";
    tmp(21516) := x"cd2d";
    tmp(21517) := x"ddae";
    tmp(21518) := x"f651";
    tmp(21519) := x"feb2";
    tmp(21520) := x"ff33";
    tmp(21521) := x"ff75";
    tmp(21522) := x"ff95";
    tmp(21523) := x"ff95";
    tmp(21524) := x"ffd6";
    tmp(21525) := x"ff74";
    tmp(21526) := x"ff33";
    tmp(21527) := x"fef1";
    tmp(21528) := x"e62f";
    tmp(21529) := x"cdad";
    tmp(21530) := x"b4ea";
    tmp(21531) := x"9c29";
    tmp(21532) := x"8387";
    tmp(21533) := x"6b05";
    tmp(21534) := x"5aa4";
    tmp(21535) := x"4a63";
    tmp(21536) := x"4223";
    tmp(21537) := x"4223";
    tmp(21538) := x"4a25";
    tmp(21539) := x"5286";
    tmp(21540) := x"5ac7";
    tmp(21541) := x"6b29";
    tmp(21542) := x"734a";
    tmp(21543) := x"836c";
    tmp(21544) := x"8bad";
    tmp(21545) := x"9c0f";
    tmp(21546) := x"a410";
    tmp(21547) := x"a451";
    tmp(21548) := x"ac51";
    tmp(21549) := x"ac71";
    tmp(21550) := x"a471";
    tmp(21551) := x"a471";
    tmp(21552) := x"9c52";
    tmp(21553) := x"9410";
    tmp(21554) := x"8bcf";
    tmp(21555) := x"7b8e";
    tmp(21556) := x"732d";
    tmp(21557) := x"f800";
    tmp(21558) := x"f800";
    tmp(21559) := x"f800";
    tmp(21560) := x"f800";
    tmp(21561) := x"f800";
    tmp(21562) := x"f800";
    tmp(21563) := x"f800";
    tmp(21564) := x"f800";
    tmp(21565) := x"f800";
    tmp(21566) := x"f800";
    tmp(21567) := x"f800";
    tmp(21568) := x"f800";
    tmp(21569) := x"f800";
    tmp(21570) := x"f800";
    tmp(21571) := x"f800";
    tmp(21572) := x"f800";
    tmp(21573) := x"f800";
    tmp(21574) := x"f800";
    tmp(21575) := x"f800";
    tmp(21576) := x"f800";
    tmp(21577) := x"f800";
    tmp(21578) := x"f800";
    tmp(21579) := x"f800";
    tmp(21580) := x"f800";
    tmp(21581) := x"f800";
    tmp(21582) := x"f800";
    tmp(21583) := x"f800";
    tmp(21584) := x"f800";
    tmp(21585) := x"f800";
    tmp(21586) := x"f800";
    tmp(21587) := x"f800";
    tmp(21588) := x"f800";
    tmp(21589) := x"f800";
    tmp(21590) := x"f800";
    tmp(21591) := x"f800";
    tmp(21592) := x"f800";
    tmp(21593) := x"f800";
    tmp(21594) := x"f800";
    tmp(21595) := x"f800";
    tmp(21596) := x"f800";
    tmp(21597) := x"0840";
    tmp(21598) := x"0840";
    tmp(21599) := x"0840";
    tmp(21600) := x"1840";
    tmp(21601) := x"fb60";
    tmp(21602) := x"eb00";
    tmp(21603) := x"eb00";
    tmp(21604) := x"fb40";
    tmp(21605) := x"f340";
    tmp(21606) := x"f340";
    tmp(21607) := x"fb60";
    tmp(21608) := x"f340";
    tmp(21609) := x"f360";
    tmp(21610) := x"fb60";
    tmp(21611) := x"fb80";
    tmp(21612) := x"fb60";
    tmp(21613) := x"fb80";
    tmp(21614) := x"fbc0";
    tmp(21615) := x"fba0";
    tmp(21616) := x"fba0";
    tmp(21617) := x"fba0";
    tmp(21618) := x"eb60";
    tmp(21619) := x"db20";
    tmp(21620) := x"db00";
    tmp(21621) := x"dac0";
    tmp(21622) := x"dac0";
    tmp(21623) := x"d2c0";
    tmp(21624) := x"caa0";
    tmp(21625) := x"ca80";
    tmp(21626) := x"cac0";
    tmp(21627) := x"cac0";
    tmp(21628) := x"dae0";
    tmp(21629) := x"dac0";
    tmp(21630) := x"eb40";
    tmp(21631) := x"f340";
    tmp(21632) := x"f340";
    tmp(21633) := x"eb40";
    tmp(21634) := x"f340";
    tmp(21635) := x"eb20";
    tmp(21636) := x"eb20";
    tmp(21637) := x"eb40";
    tmp(21638) := x"f340";
    tmp(21639) := x"fb40";
    tmp(21640) := x"fb40";
    tmp(21641) := x"fb80";
    tmp(21642) := x"f340";
    tmp(21643) := x"f340";
    tmp(21644) := x"f340";
    tmp(21645) := x"f340";
    tmp(21646) := x"fb80";
    tmp(21647) := x"fbc0";
    tmp(21648) := x"fbc0";
    tmp(21649) := x"fbc0";
    tmp(21650) := x"eb60";
    tmp(21651) := x"eb20";
    tmp(21652) := x"dac0";
    tmp(21653) := x"e2e0";
    tmp(21654) := x"eb00";
    tmp(21655) := x"eb20";
    tmp(21656) := x"eb20";
    tmp(21657) := x"eb40";
    tmp(21658) := x"db00";
    tmp(21659) := x"c2a0";
    tmp(21660) := x"c280";
    tmp(21661) := x"c2a0";
    tmp(21662) := x"cae0";
    tmp(21663) := x"d2e0";
    tmp(21664) := x"db00";
    tmp(21665) := x"db00";
    tmp(21666) := x"dae0";
    tmp(21667) := x"d2c0";
    tmp(21668) := x"d2c0";
    tmp(21669) := x"ca80";
    tmp(21670) := x"c280";
    tmp(21671) := x"ba40";
    tmp(21672) := x"ba40";
    tmp(21673) := x"c260";
    tmp(21674) := x"c280";
    tmp(21675) := x"c280";
    tmp(21676) := x"aa40";
    tmp(21677) := x"6980";
    tmp(21678) := x"28c0";
    tmp(21679) := x"0840";
    tmp(21680) := x"0020";
    tmp(21681) := x"0020";
    tmp(21682) := x"0020";
    tmp(21683) := x"0040";
    tmp(21684) := x"0840";
    tmp(21685) := x"0840";
    tmp(21686) := x"0840";
    tmp(21687) := x"0840";
    tmp(21688) := x"0860";
    tmp(21689) := x"0860";
    tmp(21690) := x"0840";
    tmp(21691) := x"0020";
    tmp(21692) := x"0000";
    tmp(21693) := x"0020";
    tmp(21694) := x"0000";
    tmp(21695) := x"0000";
    tmp(21696) := x"1040";
    tmp(21697) := x"20a0";
    tmp(21698) := x"28c0";
    tmp(21699) := x"30c0";
    tmp(21700) := x"28a0";
    tmp(21701) := x"28a0";
    tmp(21702) := x"28a0";
    tmp(21703) := x"28a0";
    tmp(21704) := x"1860";
    tmp(21705) := x"1860";
    tmp(21706) := x"30a0";
    tmp(21707) := x"5120";
    tmp(21708) := x"6960";
    tmp(21709) := x"81a0";
    tmp(21710) := x"79a0";
    tmp(21711) := x"6980";
    tmp(21712) := x"6980";
    tmp(21713) := x"79a0";
    tmp(21714) := x"8200";
    tmp(21715) := x"28c0";
    tmp(21716) := x"1060";
    tmp(21717) := x"2900";
    tmp(21718) := x"18a0";
    tmp(21719) := x"0840";
    tmp(21720) := x"3164";
    tmp(21721) := x"5a47";
    tmp(21722) := x"3984";
    tmp(21723) := x"2962";
    tmp(21724) := x"08a0";
    tmp(21725) := x"0880";
    tmp(21726) := x"0060";
    tmp(21727) := x"0060";
    tmp(21728) := x"08a0";
    tmp(21729) := x"08c0";
    tmp(21730) := x"08a0";
    tmp(21731) := x"08a0";
    tmp(21732) := x"0880";
    tmp(21733) := x"08c0";
    tmp(21734) := x"08c0";
    tmp(21735) := x"08c0";
    tmp(21736) := x"0900";
    tmp(21737) := x"1161";
    tmp(21738) := x"0921";
    tmp(21739) := x"1182";
    tmp(21740) := x"11a2";
    tmp(21741) := x"11c1";
    tmp(21742) := x"22c4";
    tmp(21743) := x"2347";
    tmp(21744) := x"2ae4";
    tmp(21745) := x"2202";
    tmp(21746) := x"1961";
    tmp(21747) := x"1941";
    tmp(21748) := x"2181";
    tmp(21749) := x"29a2";
    tmp(21750) := x"3a02";
    tmp(21751) := x"4a63";
    tmp(21752) := x"62c4";
    tmp(21753) := x"7b46";
    tmp(21754) := x"93e8";
    tmp(21755) := x"ac6a";
    tmp(21756) := x"c4ec";
    tmp(21757) := x"d58d";
    tmp(21758) := x"f630";
    tmp(21759) := x"fe71";
    tmp(21760) := x"ff13";
    tmp(21761) := x"ffb6";
    tmp(21762) := x"ff96";
    tmp(21763) := x"fff7";
    tmp(21764) := x"fff7";
    tmp(21765) := x"ffd6";
    tmp(21766) := x"ffb6";
    tmp(21767) := x"ff94";
    tmp(21768) := x"ff53";
    tmp(21769) := x"ee90";
    tmp(21770) := x"dded";
    tmp(21771) := x"bceb";
    tmp(21772) := x"a469";
    tmp(21773) := x"8ba7";
    tmp(21774) := x"7325";
    tmp(21775) := x"62c4";
    tmp(21776) := x"5264";
    tmp(21777) := x"4244";
    tmp(21778) := x"4224";
    tmp(21779) := x"52a6";
    tmp(21780) := x"5ac7";
    tmp(21781) := x"6b29";
    tmp(21782) := x"734a";
    tmp(21783) := x"838d";
    tmp(21784) := x"8bce";
    tmp(21785) := x"940f";
    tmp(21786) := x"a451";
    tmp(21787) := x"ac52";
    tmp(21788) := x"ac92";
    tmp(21789) := x"ac92";
    tmp(21790) := x"ac72";
    tmp(21791) := x"a472";
    tmp(21792) := x"a472";
    tmp(21793) := x"9c11";
    tmp(21794) := x"93f0";
    tmp(21795) := x"7b6e";
    tmp(21796) := x"734d";
    tmp(21797) := x"f800";
    tmp(21798) := x"f800";
    tmp(21799) := x"f800";
    tmp(21800) := x"f800";
    tmp(21801) := x"f800";
    tmp(21802) := x"f800";
    tmp(21803) := x"f800";
    tmp(21804) := x"f800";
    tmp(21805) := x"f800";
    tmp(21806) := x"f800";
    tmp(21807) := x"f800";
    tmp(21808) := x"f800";
    tmp(21809) := x"f800";
    tmp(21810) := x"f800";
    tmp(21811) := x"f800";
    tmp(21812) := x"f800";
    tmp(21813) := x"f800";
    tmp(21814) := x"f800";
    tmp(21815) := x"f800";
    tmp(21816) := x"f800";
    tmp(21817) := x"f800";
    tmp(21818) := x"f800";
    tmp(21819) := x"f800";
    tmp(21820) := x"f800";
    tmp(21821) := x"f800";
    tmp(21822) := x"f800";
    tmp(21823) := x"f800";
    tmp(21824) := x"f800";
    tmp(21825) := x"f800";
    tmp(21826) := x"f800";
    tmp(21827) := x"f800";
    tmp(21828) := x"f800";
    tmp(21829) := x"f800";
    tmp(21830) := x"f800";
    tmp(21831) := x"f800";
    tmp(21832) := x"f800";
    tmp(21833) := x"f800";
    tmp(21834) := x"f800";
    tmp(21835) := x"f800";
    tmp(21836) := x"f800";
    tmp(21837) := x"0840";
    tmp(21838) := x"0840";
    tmp(21839) := x"0840";
    tmp(21840) := x"1840";
    tmp(21841) := x"fb60";
    tmp(21842) := x"eb00";
    tmp(21843) := x"eb00";
    tmp(21844) := x"eae0";
    tmp(21845) := x"f340";
    tmp(21846) := x"f340";
    tmp(21847) := x"f340";
    tmp(21848) := x"f320";
    tmp(21849) := x"f320";
    tmp(21850) := x"f340";
    tmp(21851) := x"fb60";
    tmp(21852) := x"fb60";
    tmp(21853) := x"fb80";
    tmp(21854) := x"fb80";
    tmp(21855) := x"fbc0";
    tmp(21856) := x"fbe0";
    tmp(21857) := x"fc20";
    tmp(21858) := x"fc00";
    tmp(21859) := x"f360";
    tmp(21860) := x"eb20";
    tmp(21861) := x"e2e0";
    tmp(21862) := x"e2e0";
    tmp(21863) := x"e2e0";
    tmp(21864) := x"d2c0";
    tmp(21865) := x"d2c0";
    tmp(21866) := x"caa0";
    tmp(21867) := x"dac0";
    tmp(21868) := x"d2c0";
    tmp(21869) := x"dac0";
    tmp(21870) := x"dae0";
    tmp(21871) := x"f340";
    tmp(21872) := x"eb20";
    tmp(21873) := x"f340";
    tmp(21874) := x"eb20";
    tmp(21875) := x"eb20";
    tmp(21876) := x"eb00";
    tmp(21877) := x"eb20";
    tmp(21878) := x"f340";
    tmp(21879) := x"fb40";
    tmp(21880) := x"fb40";
    tmp(21881) := x"fb80";
    tmp(21882) := x"fb60";
    tmp(21883) := x"f340";
    tmp(21884) := x"f340";
    tmp(21885) := x"f340";
    tmp(21886) := x"f380";
    tmp(21887) := x"fba0";
    tmp(21888) := x"fbc0";
    tmp(21889) := x"fba0";
    tmp(21890) := x"fb80";
    tmp(21891) := x"f340";
    tmp(21892) := x"f340";
    tmp(21893) := x"f320";
    tmp(21894) := x"f320";
    tmp(21895) := x"f340";
    tmp(21896) := x"eb40";
    tmp(21897) := x"eb40";
    tmp(21898) := x"dae0";
    tmp(21899) := x"c280";
    tmp(21900) := x"c260";
    tmp(21901) := x"caa0";
    tmp(21902) := x"d2c0";
    tmp(21903) := x"d2c0";
    tmp(21904) := x"dae0";
    tmp(21905) := x"e320";
    tmp(21906) := x"db00";
    tmp(21907) := x"dae0";
    tmp(21908) := x"e2e0";
    tmp(21909) := x"e2e0";
    tmp(21910) := x"d2a0";
    tmp(21911) := x"ba60";
    tmp(21912) := x"c260";
    tmp(21913) := x"ca80";
    tmp(21914) := x"ca80";
    tmp(21915) := x"ca80";
    tmp(21916) := x"ba80";
    tmp(21917) := x"91e0";
    tmp(21918) := x"5140";
    tmp(21919) := x"20a0";
    tmp(21920) := x"0840";
    tmp(21921) := x"0840";
    tmp(21922) := x"0840";
    tmp(21923) := x"0040";
    tmp(21924) := x"0840";
    tmp(21925) := x"0840";
    tmp(21926) := x"0860";
    tmp(21927) := x"1060";
    tmp(21928) := x"1880";
    tmp(21929) := x"18a0";
    tmp(21930) := x"1080";
    tmp(21931) := x"0860";
    tmp(21932) := x"0860";
    tmp(21933) := x"1060";
    tmp(21934) := x"0840";
    tmp(21935) := x"1060";
    tmp(21936) := x"28c0";
    tmp(21937) := x"30c0";
    tmp(21938) := x"38e0";
    tmp(21939) := x"38c0";
    tmp(21940) := x"38c0";
    tmp(21941) := x"4100";
    tmp(21942) := x"5100";
    tmp(21943) := x"40c0";
    tmp(21944) := x"40c0";
    tmp(21945) := x"5920";
    tmp(21946) := x"6960";
    tmp(21947) := x"7960";
    tmp(21948) := x"89a0";
    tmp(21949) := x"89c0";
    tmp(21950) := x"89c0";
    tmp(21951) := x"81a0";
    tmp(21952) := x"81a0";
    tmp(21953) := x"9a20";
    tmp(21954) := x"69a0";
    tmp(21955) := x"20a0";
    tmp(21956) := x"2900";
    tmp(21957) := x"3100";
    tmp(21958) := x"20a0";
    tmp(21959) := x"20e1";
    tmp(21960) := x"3184";
    tmp(21961) := x"2102";
    tmp(21962) := x"10a1";
    tmp(21963) := x"0880";
    tmp(21964) := x"0880";
    tmp(21965) := x"0880";
    tmp(21966) := x"0880";
    tmp(21967) := x"0880";
    tmp(21968) := x"08a0";
    tmp(21969) := x"08a0";
    tmp(21970) := x"08a0";
    tmp(21971) := x"08a0";
    tmp(21972) := x"08a0";
    tmp(21973) := x"08c0";
    tmp(21974) := x"0900";
    tmp(21975) := x"0941";
    tmp(21976) := x"0921";
    tmp(21977) := x"0962";
    tmp(21978) := x"1183";
    tmp(21979) := x"0922";
    tmp(21980) := x"11a3";
    tmp(21981) := x"1a44";
    tmp(21982) := x"2368";
    tmp(21983) := x"33c9";
    tmp(21984) := x"3284";
    tmp(21985) := x"29c2";
    tmp(21986) := x"2181";
    tmp(21987) := x"2161";
    tmp(21988) := x"2161";
    tmp(21989) := x"2981";
    tmp(21990) := x"31c2";
    tmp(21991) := x"4243";
    tmp(21992) := x"52a4";
    tmp(21993) := x"6b05";
    tmp(21994) := x"83a7";
    tmp(21995) := x"9c09";
    tmp(21996) := x"bccb";
    tmp(21997) := x"cd6d";
    tmp(21998) := x"e5ef";
    tmp(21999) := x"f671";
    tmp(22000) := x"ff13";
    tmp(22001) := x"ff75";
    tmp(22002) := x"fff7";
    tmp(22003) := x"fff7";
    tmp(22004) := x"fff9";
    tmp(22005) := x"fffa";
    tmp(22006) := x"fff8";
    tmp(22007) := x"ffd7";
    tmp(22008) := x"fff6";
    tmp(22009) := x"ff73";
    tmp(22010) := x"f6f1";
    tmp(22011) := x"e60f";
    tmp(22012) := x"c54c";
    tmp(22013) := x"a449";
    tmp(22014) := x"8ba7";
    tmp(22015) := x"7325";
    tmp(22016) := x"5ac5";
    tmp(22017) := x"5284";
    tmp(22018) := x"4a65";
    tmp(22019) := x"5286";
    tmp(22020) := x"5ac7";
    tmp(22021) := x"6b49";
    tmp(22022) := x"736a";
    tmp(22023) := x"83cc";
    tmp(22024) := x"8bee";
    tmp(22025) := x"940f";
    tmp(22026) := x"a451";
    tmp(22027) := x"ac72";
    tmp(22028) := x"b4b3";
    tmp(22029) := x"ac93";
    tmp(22030) := x"b4b3";
    tmp(22031) := x"ac72";
    tmp(22032) := x"a452";
    tmp(22033) := x"a452";
    tmp(22034) := x"9410";
    tmp(22035) := x"838e";
    tmp(22036) := x"7b8e";
    tmp(22037) := x"f800";
    tmp(22038) := x"f800";
    tmp(22039) := x"f800";
    tmp(22040) := x"f800";
    tmp(22041) := x"f800";
    tmp(22042) := x"f800";
    tmp(22043) := x"f800";
    tmp(22044) := x"f800";
    tmp(22045) := x"f800";
    tmp(22046) := x"f800";
    tmp(22047) := x"f800";
    tmp(22048) := x"f800";
    tmp(22049) := x"f800";
    tmp(22050) := x"f800";
    tmp(22051) := x"f800";
    tmp(22052) := x"f800";
    tmp(22053) := x"f800";
    tmp(22054) := x"f800";
    tmp(22055) := x"f800";
    tmp(22056) := x"f800";
    tmp(22057) := x"f800";
    tmp(22058) := x"f800";
    tmp(22059) := x"f800";
    tmp(22060) := x"f800";
    tmp(22061) := x"f800";
    tmp(22062) := x"f800";
    tmp(22063) := x"f800";
    tmp(22064) := x"f800";
    tmp(22065) := x"f800";
    tmp(22066) := x"f800";
    tmp(22067) := x"f800";
    tmp(22068) := x"f800";
    tmp(22069) := x"f800";
    tmp(22070) := x"f800";
    tmp(22071) := x"f800";
    tmp(22072) := x"f800";
    tmp(22073) := x"f800";
    tmp(22074) := x"f800";
    tmp(22075) := x"f800";
    tmp(22076) := x"f800";
    tmp(22077) := x"0840";
    tmp(22078) := x"0840";
    tmp(22079) := x"0840";
    tmp(22080) := x"1840";
    tmp(22081) := x"fb40";
    tmp(22082) := x"eae0";
    tmp(22083) := x"eae0";
    tmp(22084) := x"eac0";
    tmp(22085) := x"fb40";
    tmp(22086) := x"fb40";
    tmp(22087) := x"fb40";
    tmp(22088) := x"fb40";
    tmp(22089) := x"fb40";
    tmp(22090) := x"fb40";
    tmp(22091) := x"fb60";
    tmp(22092) := x"f360";
    tmp(22093) := x"fb80";
    tmp(22094) := x"fb80";
    tmp(22095) := x"fbc0";
    tmp(22096) := x"fc40";
    tmp(22097) := x"fc00";
    tmp(22098) := x"fbe0";
    tmp(22099) := x"f340";
    tmp(22100) := x"eb00";
    tmp(22101) := x"eb00";
    tmp(22102) := x"f320";
    tmp(22103) := x"eb20";
    tmp(22104) := x"d2a0";
    tmp(22105) := x"d2c0";
    tmp(22106) := x"d2a0";
    tmp(22107) := x"ca80";
    tmp(22108) := x"dac0";
    tmp(22109) := x"dac0";
    tmp(22110) := x"dae0";
    tmp(22111) := x"eb20";
    tmp(22112) := x"eb20";
    tmp(22113) := x"f340";
    tmp(22114) := x"f340";
    tmp(22115) := x"f340";
    tmp(22116) := x"eb00";
    tmp(22117) := x"eb20";
    tmp(22118) := x"f340";
    tmp(22119) := x"fb40";
    tmp(22120) := x"fb60";
    tmp(22121) := x"fb40";
    tmp(22122) := x"f360";
    tmp(22123) := x"f340";
    tmp(22124) := x"f320";
    tmp(22125) := x"fb40";
    tmp(22126) := x"fb80";
    tmp(22127) := x"fbc0";
    tmp(22128) := x"fbc0";
    tmp(22129) := x"fba0";
    tmp(22130) := x"fb60";
    tmp(22131) := x"f340";
    tmp(22132) := x"fb40";
    tmp(22133) := x"fb60";
    tmp(22134) := x"fb60";
    tmp(22135) := x"fb80";
    tmp(22136) := x"f360";
    tmp(22137) := x"eb40";
    tmp(22138) := x"db00";
    tmp(22139) := x"d2c0";
    tmp(22140) := x"d2a0";
    tmp(22141) := x"d2c0";
    tmp(22142) := x"d2a0";
    tmp(22143) := x"e2e0";
    tmp(22144) := x"e2e0";
    tmp(22145) := x"eb00";
    tmp(22146) := x"eb20";
    tmp(22147) := x"eb00";
    tmp(22148) := x"eb00";
    tmp(22149) := x"eb00";
    tmp(22150) := x"dae0";
    tmp(22151) := x"ca80";
    tmp(22152) := x"ca80";
    tmp(22153) := x"ca80";
    tmp(22154) := x"c260";
    tmp(22155) := x"d2c0";
    tmp(22156) := x"c280";
    tmp(22157) := x"aa40";
    tmp(22158) := x"79c0";
    tmp(22159) := x"4920";
    tmp(22160) := x"28c0";
    tmp(22161) := x"1880";
    tmp(22162) := x"0860";
    tmp(22163) := x"0840";
    tmp(22164) := x"0840";
    tmp(22165) := x"0860";
    tmp(22166) := x"1080";
    tmp(22167) := x"1080";
    tmp(22168) := x"28e0";
    tmp(22169) := x"20c0";
    tmp(22170) := x"18a0";
    tmp(22171) := x"20c0";
    tmp(22172) := x"3920";
    tmp(22173) := x"3900";
    tmp(22174) := x"30e0";
    tmp(22175) := x"3900";
    tmp(22176) := x"30e0";
    tmp(22177) := x"4100";
    tmp(22178) := x"4920";
    tmp(22179) := x"5120";
    tmp(22180) := x"5120";
    tmp(22181) := x"5920";
    tmp(22182) := x"6120";
    tmp(22183) := x"5900";
    tmp(22184) := x"6960";
    tmp(22185) := x"7980";
    tmp(22186) := x"7980";
    tmp(22187) := x"89c0";
    tmp(22188) := x"9a00";
    tmp(22189) := x"99e0";
    tmp(22190) := x"91c0";
    tmp(22191) := x"91e0";
    tmp(22192) := x"aa40";
    tmp(22193) := x"9a00";
    tmp(22194) := x"5120";
    tmp(22195) := x"4120";
    tmp(22196) := x"4960";
    tmp(22197) := x"3920";
    tmp(22198) := x"20c0";
    tmp(22199) := x"10a0";
    tmp(22200) := x"10c1";
    tmp(22201) := x"08a0";
    tmp(22202) := x"08a0";
    tmp(22203) := x"08a0";
    tmp(22204) := x"0880";
    tmp(22205) := x"0880";
    tmp(22206) := x"08a1";
    tmp(22207) := x"08a1";
    tmp(22208) := x"08a1";
    tmp(22209) := x"08a0";
    tmp(22210) := x"08a0";
    tmp(22211) := x"08a1";
    tmp(22212) := x"08c1";
    tmp(22213) := x"0901";
    tmp(22214) := x"0961";
    tmp(22215) := x"11a3";
    tmp(22216) := x"11a4";
    tmp(22217) := x"1205";
    tmp(22218) := x"1206";
    tmp(22219) := x"1163";
    tmp(22220) := x"1204";
    tmp(22221) := x"1ac6";
    tmp(22222) := x"33aa";
    tmp(22223) := x"4347";
    tmp(22224) := x"4264";
    tmp(22225) := x"3203";
    tmp(22226) := x"29c2";
    tmp(22227) := x"2181";
    tmp(22228) := x"2161";
    tmp(22229) := x"2161";
    tmp(22230) := x"29a1";
    tmp(22231) := x"31e2";
    tmp(22232) := x"4a63";
    tmp(22233) := x"5ac4";
    tmp(22234) := x"7345";
    tmp(22235) := x"93e7";
    tmp(22236) := x"ac8a";
    tmp(22237) := x"c52b";
    tmp(22238) := x"ddae";
    tmp(22239) := x"ee50";
    tmp(22240) := x"feb2";
    tmp(22241) := x"ff54";
    tmp(22242) := x"ffd7";
    tmp(22243) := x"fff8";
    tmp(22244) := x"fff9";
    tmp(22245) := x"fffa";
    tmp(22246) := x"fffb";
    tmp(22247) := x"fff9";
    tmp(22248) := x"fff8";
    tmp(22249) := x"fff6";
    tmp(22250) := x"ff94";
    tmp(22251) := x"ff12";
    tmp(22252) := x"e630";
    tmp(22253) := x"c52c";
    tmp(22254) := x"a449";
    tmp(22255) := x"8bc7";
    tmp(22256) := x"6b26";
    tmp(22257) := x"62e5";
    tmp(22258) := x"5aa5";
    tmp(22259) := x"5ac6";
    tmp(22260) := x"5ae7";
    tmp(22261) := x"6b49";
    tmp(22262) := x"736a";
    tmp(22263) := x"7bcc";
    tmp(22264) := x"8bce";
    tmp(22265) := x"940f";
    tmp(22266) := x"9c51";
    tmp(22267) := x"a472";
    tmp(22268) := x"b4b3";
    tmp(22269) := x"b4d3";
    tmp(22270) := x"b4b2";
    tmp(22271) := x"ac72";
    tmp(22272) := x"a472";
    tmp(22273) := x"9c32";
    tmp(22274) := x"9c10";
    tmp(22275) := x"8baf";
    tmp(22276) := x"838f";
    tmp(22277) := x"f800";
    tmp(22278) := x"f800";
    tmp(22279) := x"f800";
    tmp(22280) := x"f800";
    tmp(22281) := x"f800";
    tmp(22282) := x"f800";
    tmp(22283) := x"f800";
    tmp(22284) := x"f800";
    tmp(22285) := x"f800";
    tmp(22286) := x"f800";
    tmp(22287) := x"f800";
    tmp(22288) := x"f800";
    tmp(22289) := x"f800";
    tmp(22290) := x"f800";
    tmp(22291) := x"f800";
    tmp(22292) := x"f800";
    tmp(22293) := x"f800";
    tmp(22294) := x"f800";
    tmp(22295) := x"f800";
    tmp(22296) := x"f800";
    tmp(22297) := x"f800";
    tmp(22298) := x"f800";
    tmp(22299) := x"f800";
    tmp(22300) := x"f800";
    tmp(22301) := x"f800";
    tmp(22302) := x"f800";
    tmp(22303) := x"f800";
    tmp(22304) := x"f800";
    tmp(22305) := x"f800";
    tmp(22306) := x"f800";
    tmp(22307) := x"f800";
    tmp(22308) := x"f800";
    tmp(22309) := x"f800";
    tmp(22310) := x"f800";
    tmp(22311) := x"f800";
    tmp(22312) := x"f800";
    tmp(22313) := x"f800";
    tmp(22314) := x"f800";
    tmp(22315) := x"f800";
    tmp(22316) := x"f800";
    tmp(22317) := x"0840";
    tmp(22318) := x"0840";
    tmp(22319) := x"0840";
    tmp(22320) := x"1840";
    tmp(22321) := x"f320";
    tmp(22322) := x"dac0";
    tmp(22323) := x"eae0";
    tmp(22324) := x"f300";
    tmp(22325) := x"fb40";
    tmp(22326) := x"fb60";
    tmp(22327) := x"fb40";
    tmp(22328) := x"fb40";
    tmp(22329) := x"fb40";
    tmp(22330) := x"fb40";
    tmp(22331) := x"fb60";
    tmp(22332) := x"fb60";
    tmp(22333) := x"fb80";
    tmp(22334) := x"fb80";
    tmp(22335) := x"fbc0";
    tmp(22336) := x"fbe0";
    tmp(22337) := x"fbc0";
    tmp(22338) := x"fb80";
    tmp(22339) := x"fb20";
    tmp(22340) := x"f320";
    tmp(22341) := x"f320";
    tmp(22342) := x"f320";
    tmp(22343) := x"eb20";
    tmp(22344) := x"dae0";
    tmp(22345) := x"caa0";
    tmp(22346) := x"ca80";
    tmp(22347) := x"ca60";
    tmp(22348) := x"daa0";
    tmp(22349) := x"e2c0";
    tmp(22350) := x"dac0";
    tmp(22351) := x"e2e0";
    tmp(22352) := x"e300";
    tmp(22353) := x"eb40";
    tmp(22354) := x"fb60";
    tmp(22355) := x"f340";
    tmp(22356) := x"eb40";
    tmp(22357) := x"f320";
    tmp(22358) := x"fb40";
    tmp(22359) := x"f340";
    tmp(22360) := x"fb60";
    tmp(22361) := x"fb80";
    tmp(22362) := x"f360";
    tmp(22363) := x"f340";
    tmp(22364) := x"eb00";
    tmp(22365) := x"fb40";
    tmp(22366) := x"fb60";
    tmp(22367) := x"fba0";
    tmp(22368) := x"fbc0";
    tmp(22369) := x"fba0";
    tmp(22370) := x"fba0";
    tmp(22371) := x"fb80";
    tmp(22372) := x"fb60";
    tmp(22373) := x"fb80";
    tmp(22374) := x"fba0";
    tmp(22375) := x"fb80";
    tmp(22376) := x"fbc0";
    tmp(22377) := x"f380";
    tmp(22378) := x"eb40";
    tmp(22379) := x"e2e0";
    tmp(22380) := x"dac0";
    tmp(22381) := x"dac0";
    tmp(22382) := x"ca80";
    tmp(22383) := x"dac0";
    tmp(22384) := x"eae0";
    tmp(22385) := x"eb00";
    tmp(22386) := x"f340";
    tmp(22387) := x"fb60";
    tmp(22388) := x"fb60";
    tmp(22389) := x"fb40";
    tmp(22390) := x"eb20";
    tmp(22391) := x"e300";
    tmp(22392) := x"d280";
    tmp(22393) := x"d280";
    tmp(22394) := x"ca80";
    tmp(22395) := x"d280";
    tmp(22396) := x"ca80";
    tmp(22397) := x"ba60";
    tmp(22398) := x"aa40";
    tmp(22399) := x"9200";
    tmp(22400) := x"69a0";
    tmp(22401) := x"38e0";
    tmp(22402) := x"18a0";
    tmp(22403) := x"1080";
    tmp(22404) := x"1080";
    tmp(22405) := x"1080";
    tmp(22406) := x"18a0";
    tmp(22407) := x"20a0";
    tmp(22408) := x"30e0";
    tmp(22409) := x"30e0";
    tmp(22410) := x"3920";
    tmp(22411) := x"5160";
    tmp(22412) := x"71c0";
    tmp(22413) := x"5960";
    tmp(22414) := x"5960";
    tmp(22415) := x"5940";
    tmp(22416) := x"5140";
    tmp(22417) := x"6180";
    tmp(22418) := x"6980";
    tmp(22419) := x"6980";
    tmp(22420) := x"6960";
    tmp(22421) := x"6940";
    tmp(22422) := x"7140";
    tmp(22423) := x"7960";
    tmp(22424) := x"81a0";
    tmp(22425) := x"89a0";
    tmp(22426) := x"99e0";
    tmp(22427) := x"aa20";
    tmp(22428) := x"aa00";
    tmp(22429) := x"99e0";
    tmp(22430) := x"a200";
    tmp(22431) := x"aa40";
    tmp(22432) := x"b240";
    tmp(22433) := x"91e0";
    tmp(22434) := x"6980";
    tmp(22435) := x"61a0";
    tmp(22436) := x"4140";
    tmp(22437) := x"20e0";
    tmp(22438) := x"1080";
    tmp(22439) := x"08a0";
    tmp(22440) := x"0880";
    tmp(22441) := x"08a0";
    tmp(22442) := x"08a0";
    tmp(22443) := x"08a0";
    tmp(22444) := x"08a1";
    tmp(22445) := x"08a1";
    tmp(22446) := x"08a1";
    tmp(22447) := x"08a1";
    tmp(22448) := x"08c1";
    tmp(22449) := x"08c1";
    tmp(22450) := x"08e1";
    tmp(22451) := x"08c1";
    tmp(22452) := x"0901";
    tmp(22453) := x"0922";
    tmp(22454) := x"0942";
    tmp(22455) := x"11a3";
    tmp(22456) := x"1a66";
    tmp(22457) := x"1aa8";
    tmp(22458) := x"1206";
    tmp(22459) := x"1a46";
    tmp(22460) := x"22c8";
    tmp(22461) := x"334a";
    tmp(22462) := x"53a9";
    tmp(22463) := x"5306";
    tmp(22464) := x"4a84";
    tmp(22465) := x"4264";
    tmp(22466) := x"3a23";
    tmp(22467) := x"31e2";
    tmp(22468) := x"29a1";
    tmp(22469) := x"2181";
    tmp(22470) := x"2181";
    tmp(22471) := x"29a1";
    tmp(22472) := x"3a02";
    tmp(22473) := x"4a83";
    tmp(22474) := x"6b04";
    tmp(22475) := x"8386";
    tmp(22476) := x"9c28";
    tmp(22477) := x"b4ca";
    tmp(22478) := x"cd4c";
    tmp(22479) := x"edef";
    tmp(22480) := x"fe91";
    tmp(22481) := x"ff34";
    tmp(22482) := x"ffb6";
    tmp(22483) := x"fff9";
    tmp(22484) := x"fffb";
    tmp(22485) := x"fffc";
    tmp(22486) := x"fffc";
    tmp(22487) := x"fffc";
    tmp(22488) := x"fffa";
    tmp(22489) := x"fff8";
    tmp(22490) := x"fff7";
    tmp(22491) := x"ff95";
    tmp(22492) := x"fef2";
    tmp(22493) := x"ee0f";
    tmp(22494) := x"c52c";
    tmp(22495) := x"9c49";
    tmp(22496) := x"83a7";
    tmp(22497) := x"7346";
    tmp(22498) := x"62c6";
    tmp(22499) := x"5ac6";
    tmp(22500) := x"62e8";
    tmp(22501) := x"6b4a";
    tmp(22502) := x"736b";
    tmp(22503) := x"7bcd";
    tmp(22504) := x"8c0e";
    tmp(22505) := x"9430";
    tmp(22506) := x"9c51";
    tmp(22507) := x"a472";
    tmp(22508) := x"ac93";
    tmp(22509) := x"b4d3";
    tmp(22510) := x"bcd3";
    tmp(22511) := x"b493";
    tmp(22512) := x"ac93";
    tmp(22513) := x"ac52";
    tmp(22514) := x"a452";
    tmp(22515) := x"93d0";
    tmp(22516) := x"8baf";
    tmp(22517) := x"f800";
    tmp(22518) := x"f800";
    tmp(22519) := x"f800";
    tmp(22520) := x"f800";
    tmp(22521) := x"f800";
    tmp(22522) := x"f800";
    tmp(22523) := x"f800";
    tmp(22524) := x"f800";
    tmp(22525) := x"f800";
    tmp(22526) := x"f800";
    tmp(22527) := x"f800";
    tmp(22528) := x"f800";
    tmp(22529) := x"f800";
    tmp(22530) := x"f800";
    tmp(22531) := x"f800";
    tmp(22532) := x"f800";
    tmp(22533) := x"f800";
    tmp(22534) := x"f800";
    tmp(22535) := x"f800";
    tmp(22536) := x"f800";
    tmp(22537) := x"f800";
    tmp(22538) := x"f800";
    tmp(22539) := x"f800";
    tmp(22540) := x"f800";
    tmp(22541) := x"f800";
    tmp(22542) := x"f800";
    tmp(22543) := x"f800";
    tmp(22544) := x"f800";
    tmp(22545) := x"f800";
    tmp(22546) := x"f800";
    tmp(22547) := x"f800";
    tmp(22548) := x"f800";
    tmp(22549) := x"f800";
    tmp(22550) := x"f800";
    tmp(22551) := x"f800";
    tmp(22552) := x"f800";
    tmp(22553) := x"f800";
    tmp(22554) := x"f800";
    tmp(22555) := x"f800";
    tmp(22556) := x"f800";
    tmp(22557) := x"0840";
    tmp(22558) := x"0840";
    tmp(22559) := x"0840";
    tmp(22560) := x"1840";
    tmp(22561) := x"f320";
    tmp(22562) := x"e2e0";
    tmp(22563) := x"eb00";
    tmp(22564) := x"f300";
    tmp(22565) := x"f320";
    tmp(22566) := x"fb40";
    tmp(22567) := x"fb40";
    tmp(22568) := x"fb20";
    tmp(22569) := x"fb40";
    tmp(22570) := x"fb40";
    tmp(22571) := x"fb40";
    tmp(22572) := x"fb40";
    tmp(22573) := x"fb60";
    tmp(22574) := x"fb80";
    tmp(22575) := x"fba0";
    tmp(22576) := x"fbe0";
    tmp(22577) := x"fbc0";
    tmp(22578) := x"fb80";
    tmp(22579) := x"fb20";
    tmp(22580) := x"f300";
    tmp(22581) := x"eb00";
    tmp(22582) := x"eb00";
    tmp(22583) := x"eb20";
    tmp(22584) := x"f320";
    tmp(22585) := x"dae0";
    tmp(22586) := x"d2a0";
    tmp(22587) := x"daa0";
    tmp(22588) := x"da80";
    tmp(22589) := x"daa0";
    tmp(22590) := x"eac0";
    tmp(22591) := x"e2e0";
    tmp(22592) := x"e2e0";
    tmp(22593) := x"f340";
    tmp(22594) := x"eb20";
    tmp(22595) := x"f320";
    tmp(22596) := x"fb40";
    tmp(22597) := x"f340";
    tmp(22598) := x"f340";
    tmp(22599) := x"fb40";
    tmp(22600) := x"fb40";
    tmp(22601) := x"f360";
    tmp(22602) := x"f340";
    tmp(22603) := x"f340";
    tmp(22604) := x"f300";
    tmp(22605) := x"fb40";
    tmp(22606) := x"fb60";
    tmp(22607) := x"fba0";
    tmp(22608) := x"fb80";
    tmp(22609) := x"fba0";
    tmp(22610) := x"fba0";
    tmp(22611) := x"fba0";
    tmp(22612) := x"fba0";
    tmp(22613) := x"fb80";
    tmp(22614) := x"fba0";
    tmp(22615) := x"fba0";
    tmp(22616) := x"fbc0";
    tmp(22617) := x"fbc0";
    tmp(22618) := x"fba0";
    tmp(22619) := x"fb40";
    tmp(22620) := x"e2e0";
    tmp(22621) := x"ca60";
    tmp(22622) := x"d280";
    tmp(22623) := x"eae0";
    tmp(22624) := x"eb00";
    tmp(22625) := x"fb40";
    tmp(22626) := x"fb40";
    tmp(22627) := x"fb80";
    tmp(22628) := x"fbc0";
    tmp(22629) := x"fb60";
    tmp(22630) := x"fb80";
    tmp(22631) := x"f340";
    tmp(22632) := x"e2e0";
    tmp(22633) := x"dac0";
    tmp(22634) := x"d2a0";
    tmp(22635) := x"ca80";
    tmp(22636) := x"ca80";
    tmp(22637) := x"ca80";
    tmp(22638) := x"c280";
    tmp(22639) := x"c280";
    tmp(22640) := x"a220";
    tmp(22641) := x"71a0";
    tmp(22642) := x"5140";
    tmp(22643) := x"4120";
    tmp(22644) := x"4120";
    tmp(22645) := x"3900";
    tmp(22646) := x"4120";
    tmp(22647) := x"4120";
    tmp(22648) := x"5980";
    tmp(22649) := x"69a0";
    tmp(22650) := x"71e0";
    tmp(22651) := x"8a20";
    tmp(22652) := x"9220";
    tmp(22653) := x"81e0";
    tmp(22654) := x"79c0";
    tmp(22655) := x"7180";
    tmp(22656) := x"79a0";
    tmp(22657) := x"89e0";
    tmp(22658) := x"79a0";
    tmp(22659) := x"7180";
    tmp(22660) := x"7160";
    tmp(22661) := x"7140";
    tmp(22662) := x"8980";
    tmp(22663) := x"91c0";
    tmp(22664) := x"8980";
    tmp(22665) := x"a1e0";
    tmp(22666) := x"ba40";
    tmp(22667) := x"b220";
    tmp(22668) := x"b200";
    tmp(22669) := x"aa00";
    tmp(22670) := x"aa20";
    tmp(22671) := x"ba60";
    tmp(22672) := x"aa40";
    tmp(22673) := x"81c0";
    tmp(22674) := x"6180";
    tmp(22675) := x"4160";
    tmp(22676) := x"1900";
    tmp(22677) := x"08c0";
    tmp(22678) := x"08a0";
    tmp(22679) := x"08a0";
    tmp(22680) := x"08c0";
    tmp(22681) := x"08c0";
    tmp(22682) := x"08c0";
    tmp(22683) := x"00a0";
    tmp(22684) := x"00a1";
    tmp(22685) := x"00a2";
    tmp(22686) := x"08c2";
    tmp(22687) := x"0902";
    tmp(22688) := x"08e2";
    tmp(22689) := x"08e1";
    tmp(22690) := x"0902";
    tmp(22691) := x"0922";
    tmp(22692) := x"0943";
    tmp(22693) := x"0923";
    tmp(22694) := x"0963";
    tmp(22695) := x"1204";
    tmp(22696) := x"1ac8";
    tmp(22697) := x"1267";
    tmp(22698) := x"1247";
    tmp(22699) := x"234b";
    tmp(22700) := x"440d";
    tmp(22701) := x"74cc";
    tmp(22702) := x"73c8";
    tmp(22703) := x"6b47";
    tmp(22704) := x"5ae5";
    tmp(22705) := x"52a4";
    tmp(22706) := x"4a64";
    tmp(22707) := x"3a23";
    tmp(22708) := x"31e2";
    tmp(22709) := x"29a2";
    tmp(22710) := x"2181";
    tmp(22711) := x"2181";
    tmp(22712) := x"31c2";
    tmp(22713) := x"4242";
    tmp(22714) := x"52a4";
    tmp(22715) := x"6b45";
    tmp(22716) := x"8bc7";
    tmp(22717) := x"a469";
    tmp(22718) := x"c50b";
    tmp(22719) := x"ddad";
    tmp(22720) := x"f670";
    tmp(22721) := x"ff12";
    tmp(22722) := x"ffb5";
    tmp(22723) := x"fff8";
    tmp(22724) := x"fffa";
    tmp(22725) := x"fffd";
    tmp(22726) := x"fffe";
    tmp(22727) := x"fffe";
    tmp(22728) := x"fffd";
    tmp(22729) := x"fffb";
    tmp(22730) := x"fffa";
    tmp(22731) := x"ffd8";
    tmp(22732) := x"ffb6";
    tmp(22733) := x"ff12";
    tmp(22734) := x"ee0f";
    tmp(22735) := x"bceb";
    tmp(22736) := x"9c49";
    tmp(22737) := x"83a7";
    tmp(22738) := x"6b27";
    tmp(22739) := x"62c7";
    tmp(22740) := x"6308";
    tmp(22741) := x"734a";
    tmp(22742) := x"7b8c";
    tmp(22743) := x"83ed";
    tmp(22744) := x"8c0e";
    tmp(22745) := x"9c50";
    tmp(22746) := x"a471";
    tmp(22747) := x"ac72";
    tmp(22748) := x"ac93";
    tmp(22749) := x"bcd3";
    tmp(22750) := x"c4f4";
    tmp(22751) := x"bcd4";
    tmp(22752) := x"b4d4";
    tmp(22753) := x"ac72";
    tmp(22754) := x"ac92";
    tmp(22755) := x"9c11";
    tmp(22756) := x"93f0";
    tmp(22757) := x"f800";
    tmp(22758) := x"f800";
    tmp(22759) := x"f800";
    tmp(22760) := x"f800";
    tmp(22761) := x"f800";
    tmp(22762) := x"f800";
    tmp(22763) := x"f800";
    tmp(22764) := x"f800";
    tmp(22765) := x"f800";
    tmp(22766) := x"f800";
    tmp(22767) := x"f800";
    tmp(22768) := x"f800";
    tmp(22769) := x"f800";
    tmp(22770) := x"f800";
    tmp(22771) := x"f800";
    tmp(22772) := x"f800";
    tmp(22773) := x"f800";
    tmp(22774) := x"f800";
    tmp(22775) := x"f800";
    tmp(22776) := x"f800";
    tmp(22777) := x"f800";
    tmp(22778) := x"f800";
    tmp(22779) := x"f800";
    tmp(22780) := x"f800";
    tmp(22781) := x"f800";
    tmp(22782) := x"f800";
    tmp(22783) := x"f800";
    tmp(22784) := x"f800";
    tmp(22785) := x"f800";
    tmp(22786) := x"f800";
    tmp(22787) := x"f800";
    tmp(22788) := x"f800";
    tmp(22789) := x"f800";
    tmp(22790) := x"f800";
    tmp(22791) := x"f800";
    tmp(22792) := x"f800";
    tmp(22793) := x"f800";
    tmp(22794) := x"f800";
    tmp(22795) := x"f800";
    tmp(22796) := x"f800";
    tmp(22797) := x"0840";
    tmp(22798) := x"0840";
    tmp(22799) := x"0840";
    tmp(22800) := x"1040";
    tmp(22801) := x"e300";
    tmp(22802) := x"dac0";
    tmp(22803) := x"eae0";
    tmp(22804) := x"f300";
    tmp(22805) := x"f300";
    tmp(22806) := x"fb20";
    tmp(22807) := x"fb20";
    tmp(22808) := x"fb00";
    tmp(22809) := x"fb20";
    tmp(22810) := x"fb20";
    tmp(22811) := x"fb20";
    tmp(22812) := x"fb40";
    tmp(22813) := x"fb40";
    tmp(22814) := x"fb60";
    tmp(22815) := x"fb80";
    tmp(22816) := x"fb80";
    tmp(22817) := x"fb80";
    tmp(22818) := x"fb40";
    tmp(22819) := x"f320";
    tmp(22820) := x"eae0";
    tmp(22821) := x"eae0";
    tmp(22822) := x"f320";
    tmp(22823) := x"f320";
    tmp(22824) := x"f340";
    tmp(22825) := x"eb20";
    tmp(22826) := x"eb00";
    tmp(22827) := x"e2e0";
    tmp(22828) := x"daa0";
    tmp(22829) := x"daa0";
    tmp(22830) := x"daa0";
    tmp(22831) := x"e2e0";
    tmp(22832) := x"f320";
    tmp(22833) := x"d2a0";
    tmp(22834) := x"ca80";
    tmp(22835) := x"eb20";
    tmp(22836) := x"f340";
    tmp(22837) := x"fb80";
    tmp(22838) := x"fb80";
    tmp(22839) := x"fb80";
    tmp(22840) := x"f360";
    tmp(22841) := x"f340";
    tmp(22842) := x"f360";
    tmp(22843) := x"eb20";
    tmp(22844) := x"f340";
    tmp(22845) := x"fb40";
    tmp(22846) := x"f340";
    tmp(22847) := x"fb60";
    tmp(22848) := x"fb80";
    tmp(22849) := x"fbc0";
    tmp(22850) := x"fbc0";
    tmp(22851) := x"fbc0";
    tmp(22852) := x"fbc0";
    tmp(22853) := x"fba0";
    tmp(22854) := x"fb80";
    tmp(22855) := x"fba0";
    tmp(22856) := x"fbe0";
    tmp(22857) := x"fbe0";
    tmp(22858) := x"fba0";
    tmp(22859) := x"fb60";
    tmp(22860) := x"eae0";
    tmp(22861) := x"da80";
    tmp(22862) := x"da80";
    tmp(22863) := x"eac0";
    tmp(22864) := x"f2e0";
    tmp(22865) := x"fb20";
    tmp(22866) := x"fb40";
    tmp(22867) := x"fb80";
    tmp(22868) := x"fba0";
    tmp(22869) := x"fc00";
    tmp(22870) := x"fbe0";
    tmp(22871) := x"fc00";
    tmp(22872) := x"eb40";
    tmp(22873) := x"d2a0";
    tmp(22874) := x"dac0";
    tmp(22875) := x"dac0";
    tmp(22876) := x"dac0";
    tmp(22877) := x"d2c0";
    tmp(22878) := x"d2a0";
    tmp(22879) := x"ca60";
    tmp(22880) := x"ca80";
    tmp(22881) := x"ba60";
    tmp(22882) := x"aa40";
    tmp(22883) := x"aa40";
    tmp(22884) := x"9a20";
    tmp(22885) := x"9200";
    tmp(22886) := x"9a20";
    tmp(22887) := x"9200";
    tmp(22888) := x"aa60";
    tmp(22889) := x"b280";
    tmp(22890) := x"9a40";
    tmp(22891) := x"b280";
    tmp(22892) := x"bac0";
    tmp(22893) := x"a220";
    tmp(22894) := x"91e0";
    tmp(22895) := x"89c0";
    tmp(22896) := x"91e0";
    tmp(22897) := x"91e0";
    tmp(22898) := x"89a0";
    tmp(22899) := x"7960";
    tmp(22900) := x"7980";
    tmp(22901) := x"89a0";
    tmp(22902) := x"91a0";
    tmp(22903) := x"91a0";
    tmp(22904) := x"99e0";
    tmp(22905) := x"a1e0";
    tmp(22906) := x"aa20";
    tmp(22907) := x"a1e0";
    tmp(22908) := x"aa00";
    tmp(22909) := x"b220";
    tmp(22910) := x"b240";
    tmp(22911) := x"b240";
    tmp(22912) := x"9200";
    tmp(22913) := x"5980";
    tmp(22914) := x"3140";
    tmp(22915) := x"10e0";
    tmp(22916) := x"08c0";
    tmp(22917) := x"08c0";
    tmp(22918) := x"08c0";
    tmp(22919) := x"08c1";
    tmp(22920) := x"08c0";
    tmp(22921) := x"08a0";
    tmp(22922) := x"08a0";
    tmp(22923) := x"00a0";
    tmp(22924) := x"08c1";
    tmp(22925) := x"08e2";
    tmp(22926) := x"08e2";
    tmp(22927) := x"08e2";
    tmp(22928) := x"08e2";
    tmp(22929) := x"0903";
    tmp(22930) := x"0923";
    tmp(22931) := x"0963";
    tmp(22932) := x"0964";
    tmp(22933) := x"0943";
    tmp(22934) := x"0984";
    tmp(22935) := x"1267";
    tmp(22936) := x"1289";
    tmp(22937) := x"1227";
    tmp(22938) := x"22c9";
    tmp(22939) := x"548e";
    tmp(22940) := x"956e";
    tmp(22941) := x"94aa";
    tmp(22942) := x"8c09";
    tmp(22943) := x"7ba8";
    tmp(22944) := x"6b47";
    tmp(22945) := x"6306";
    tmp(22946) := x"5ac5";
    tmp(22947) := x"4a84";
    tmp(22948) := x"3a23";
    tmp(22949) := x"3202";
    tmp(22950) := x"29a2";
    tmp(22951) := x"2981";
    tmp(22952) := x"29a1";
    tmp(22953) := x"31e2";
    tmp(22954) := x"4a63";
    tmp(22955) := x"62e4";
    tmp(22956) := x"7b46";
    tmp(22957) := x"93e7";
    tmp(22958) := x"acaa";
    tmp(22959) := x"cd4c";
    tmp(22960) := x"e62f";
    tmp(22961) := x"fed2";
    tmp(22962) := x"ff74";
    tmp(22963) := x"ffd7";
    tmp(22964) := x"fff8";
    tmp(22965) := x"fffc";
    tmp(22966) := x"fffe";
    tmp(22967) := x"ffff";
    tmp(22968) := x"ffff";
    tmp(22969) := x"fffe";
    tmp(22970) := x"fffd";
    tmp(22971) := x"fffb";
    tmp(22972) := x"fff8";
    tmp(22973) := x"ff95";
    tmp(22974) := x"fed2";
    tmp(22975) := x"d58d";
    tmp(22976) := x"bceb";
    tmp(22977) := x"9c69";
    tmp(22978) := x"7b68";
    tmp(22979) := x"6b08";
    tmp(22980) := x"6308";
    tmp(22981) := x"736b";
    tmp(22982) := x"83ac";
    tmp(22983) := x"8bee";
    tmp(22984) := x"8c0e";
    tmp(22985) := x"9c70";
    tmp(22986) := x"a491";
    tmp(22987) := x"a471";
    tmp(22988) := x"ac92";
    tmp(22989) := x"b4d3";
    tmp(22990) := x"bcf4";
    tmp(22991) := x"bcf5";
    tmp(22992) := x"b4d3";
    tmp(22993) := x"b4d2";
    tmp(22994) := x"a472";
    tmp(22995) := x"a472";
    tmp(22996) := x"9c12";
    tmp(22997) := x"f800";
    tmp(22998) := x"f800";
    tmp(22999) := x"f800";
    tmp(23000) := x"f800";
    tmp(23001) := x"f800";
    tmp(23002) := x"f800";
    tmp(23003) := x"f800";
    tmp(23004) := x"f800";
    tmp(23005) := x"f800";
    tmp(23006) := x"f800";
    tmp(23007) := x"f800";
    tmp(23008) := x"f800";
    tmp(23009) := x"f800";
    tmp(23010) := x"f800";
    tmp(23011) := x"f800";
    tmp(23012) := x"f800";
    tmp(23013) := x"f800";
    tmp(23014) := x"f800";
    tmp(23015) := x"f800";
    tmp(23016) := x"f800";
    tmp(23017) := x"f800";
    tmp(23018) := x"f800";
    tmp(23019) := x"f800";
    tmp(23020) := x"f800";
    tmp(23021) := x"f800";
    tmp(23022) := x"f800";
    tmp(23023) := x"f800";
    tmp(23024) := x"f800";
    tmp(23025) := x"f800";
    tmp(23026) := x"f800";
    tmp(23027) := x"f800";
    tmp(23028) := x"f800";
    tmp(23029) := x"f800";
    tmp(23030) := x"f800";
    tmp(23031) := x"f800";
    tmp(23032) := x"f800";
    tmp(23033) := x"f800";
    tmp(23034) := x"f800";
    tmp(23035) := x"f800";
    tmp(23036) := x"f800";
    tmp(23037) := x"0840";
    tmp(23038) := x"0840";
    tmp(23039) := x"0840";
    tmp(23040) := x"1040";
    tmp(23041) := x"e2e0";
    tmp(23042) := x"dac0";
    tmp(23043) := x"eae0";
    tmp(23044) := x"eb00";
    tmp(23045) := x"f300";
    tmp(23046) := x"fb20";
    tmp(23047) := x"fb00";
    tmp(23048) := x"fb20";
    tmp(23049) := x"fb00";
    tmp(23050) := x"fae0";
    tmp(23051) := x"fb00";
    tmp(23052) := x"fb20";
    tmp(23053) := x"fb20";
    tmp(23054) := x"fb40";
    tmp(23055) := x"fb40";
    tmp(23056) := x"fb60";
    tmp(23057) := x"fb60";
    tmp(23058) := x"fb40";
    tmp(23059) := x"eb00";
    tmp(23060) := x"eac0";
    tmp(23061) := x"f300";
    tmp(23062) := x"eb00";
    tmp(23063) := x"f320";
    tmp(23064) := x"fb40";
    tmp(23065) := x"fb60";
    tmp(23066) := x"f340";
    tmp(23067) := x"eb00";
    tmp(23068) := x"eae0";
    tmp(23069) := x"daa0";
    tmp(23070) := x"e2c0";
    tmp(23071) := x"dac0";
    tmp(23072) := x"ca80";
    tmp(23073) := x"ca60";
    tmp(23074) := x"e300";
    tmp(23075) := x"eb40";
    tmp(23076) := x"f340";
    tmp(23077) := x"fb60";
    tmp(23078) := x"fb60";
    tmp(23079) := x"fb60";
    tmp(23080) := x"fb60";
    tmp(23081) := x"eb40";
    tmp(23082) := x"f360";
    tmp(23083) := x"eb20";
    tmp(23084) := x"f340";
    tmp(23085) := x"eb20";
    tmp(23086) := x"eb40";
    tmp(23087) := x"f360";
    tmp(23088) := x"fb80";
    tmp(23089) := x"fba0";
    tmp(23090) := x"fbe0";
    tmp(23091) := x"fbc0";
    tmp(23092) := x"fba0";
    tmp(23093) := x"fb80";
    tmp(23094) := x"fb80";
    tmp(23095) := x"fbc0";
    tmp(23096) := x"fba0";
    tmp(23097) := x"fbe0";
    tmp(23098) := x"fc00";
    tmp(23099) := x"fb80";
    tmp(23100) := x"f320";
    tmp(23101) := x"e2c0";
    tmp(23102) := x"da80";
    tmp(23103) := x"e280";
    tmp(23104) := x"f2c0";
    tmp(23105) := x"fb00";
    tmp(23106) := x"fb60";
    tmp(23107) := x"fb40";
    tmp(23108) := x"fba0";
    tmp(23109) := x"fc00";
    tmp(23110) := x"fc80";
    tmp(23111) := x"fc40";
    tmp(23112) := x"fb80";
    tmp(23113) := x"eb00";
    tmp(23114) := x"eae0";
    tmp(23115) := x"eb00";
    tmp(23116) := x"eb00";
    tmp(23117) := x"e2e0";
    tmp(23118) := x"daa0";
    tmp(23119) := x"d280";
    tmp(23120) := x"daa0";
    tmp(23121) := x"dac0";
    tmp(23122) := x"eb00";
    tmp(23123) := x"eb20";
    tmp(23124) := x"e2e0";
    tmp(23125) := x"d2a0";
    tmp(23126) := x"c260";
    tmp(23127) := x"c280";
    tmp(23128) := x"eb20";
    tmp(23129) := x"ba80";
    tmp(23130) := x"c2c0";
    tmp(23131) := x"db20";
    tmp(23132) := x"dac0";
    tmp(23133) := x"ba40";
    tmp(23134) := x"a1e0";
    tmp(23135) := x"a200";
    tmp(23136) := x"aa20";
    tmp(23137) := x"99e0";
    tmp(23138) := x"89a0";
    tmp(23139) := x"8180";
    tmp(23140) := x"89a0";
    tmp(23141) := x"91c0";
    tmp(23142) := x"99c0";
    tmp(23143) := x"aa00";
    tmp(23144) := x"99c0";
    tmp(23145) := x"99c0";
    tmp(23146) := x"91c0";
    tmp(23147) := x"99e0";
    tmp(23148) := x"aa20";
    tmp(23149) := x"aa20";
    tmp(23150) := x"aa40";
    tmp(23151) := x"aa60";
    tmp(23152) := x"71e0";
    tmp(23153) := x"2920";
    tmp(23154) := x"10c0";
    tmp(23155) := x"08c0";
    tmp(23156) := x"08c0";
    tmp(23157) := x"08c1";
    tmp(23158) := x"08e1";
    tmp(23159) := x"08c1";
    tmp(23160) := x"08c1";
    tmp(23161) := x"08c0";
    tmp(23162) := x"08c1";
    tmp(23163) := x"0901";
    tmp(23164) := x"0923";
    tmp(23165) := x"08c2";
    tmp(23166) := x"08e2";
    tmp(23167) := x"0923";
    tmp(23168) := x"0904";
    tmp(23169) := x"0924";
    tmp(23170) := x"0924";
    tmp(23171) := x"0965";
    tmp(23172) := x"0965";
    tmp(23173) := x"11a6";
    tmp(23174) := x"1207";
    tmp(23175) := x"1acb";
    tmp(23176) := x"1249";
    tmp(23177) := x"2289";
    tmp(23178) := x"6ccf";
    tmp(23179) := x"a5ae";
    tmp(23180) := x"b52c";
    tmp(23181) := x"aceb";
    tmp(23182) := x"9c8a";
    tmp(23183) := x"9449";
    tmp(23184) := x"83c8";
    tmp(23185) := x"7367";
    tmp(23186) := x"6b46";
    tmp(23187) := x"5ae5";
    tmp(23188) := x"5284";
    tmp(23189) := x"4243";
    tmp(23190) := x"3a03";
    tmp(23191) := x"31c2";
    tmp(23192) := x"29a2";
    tmp(23193) := x"31a2";
    tmp(23194) := x"3a22";
    tmp(23195) := x"5283";
    tmp(23196) := x"6ae5";
    tmp(23197) := x"83a6";
    tmp(23198) := x"9c68";
    tmp(23199) := x"b4ea";
    tmp(23200) := x"d5ad";
    tmp(23201) := x"f670";
    tmp(23202) := x"ff12";
    tmp(23203) := x"ffb5";
    tmp(23204) := x"fff8";
    tmp(23205) := x"fffc";
    tmp(23206) := x"ffff";
    tmp(23207) := x"ffff";
    tmp(23208) := x"ffff";
    tmp(23209) := x"ffff";
    tmp(23210) := x"ffff";
    tmp(23211) := x"fffe";
    tmp(23212) := x"fffc";
    tmp(23213) := x"fff8";
    tmp(23214) := x"ff34";
    tmp(23215) := x"ee0f";
    tmp(23216) := x"d5ad";
    tmp(23217) := x"b4cb";
    tmp(23218) := x"8bca";
    tmp(23219) := x"6b28";
    tmp(23220) := x"6309";
    tmp(23221) := x"736b";
    tmp(23222) := x"83cd";
    tmp(23223) := x"8bcd";
    tmp(23224) := x"9450";
    tmp(23225) := x"9c71";
    tmp(23226) := x"a492";
    tmp(23227) := x"a4b2";
    tmp(23228) := x"acb2";
    tmp(23229) := x"b4d3";
    tmp(23230) := x"c535";
    tmp(23231) := x"bcf5";
    tmp(23232) := x"bd14";
    tmp(23233) := x"b4d3";
    tmp(23234) := x"acb3";
    tmp(23235) := x"a472";
    tmp(23236) := x"a453";
    tmp(23237) := x"f800";
    tmp(23238) := x"f800";
    tmp(23239) := x"f800";
    tmp(23240) := x"f800";
    tmp(23241) := x"f800";
    tmp(23242) := x"f800";
    tmp(23243) := x"f800";
    tmp(23244) := x"f800";
    tmp(23245) := x"f800";
    tmp(23246) := x"f800";
    tmp(23247) := x"f800";
    tmp(23248) := x"f800";
    tmp(23249) := x"f800";
    tmp(23250) := x"f800";
    tmp(23251) := x"f800";
    tmp(23252) := x"f800";
    tmp(23253) := x"f800";
    tmp(23254) := x"f800";
    tmp(23255) := x"f800";
    tmp(23256) := x"f800";
    tmp(23257) := x"f800";
    tmp(23258) := x"f800";
    tmp(23259) := x"f800";
    tmp(23260) := x"f800";
    tmp(23261) := x"f800";
    tmp(23262) := x"f800";
    tmp(23263) := x"f800";
    tmp(23264) := x"f800";
    tmp(23265) := x"f800";
    tmp(23266) := x"f800";
    tmp(23267) := x"f800";
    tmp(23268) := x"f800";
    tmp(23269) := x"f800";
    tmp(23270) := x"f800";
    tmp(23271) := x"f800";
    tmp(23272) := x"f800";
    tmp(23273) := x"f800";
    tmp(23274) := x"f800";
    tmp(23275) := x"f800";
    tmp(23276) := x"f800";
    tmp(23277) := x"0840";
    tmp(23278) := x"0840";
    tmp(23279) := x"0840";
    tmp(23280) := x"1040";
    tmp(23281) := x"eb40";
    tmp(23282) := x"dae0";
    tmp(23283) := x"eb20";
    tmp(23284) := x"eb20";
    tmp(23285) := x"fb40";
    tmp(23286) := x"fb40";
    tmp(23287) := x"fb40";
    tmp(23288) := x"fb40";
    tmp(23289) := x"fb40";
    tmp(23290) := x"fb00";
    tmp(23291) := x"fb00";
    tmp(23292) := x"fb00";
    tmp(23293) := x"fb20";
    tmp(23294) := x"fb20";
    tmp(23295) := x"fb60";
    tmp(23296) := x"fb60";
    tmp(23297) := x"fb40";
    tmp(23298) := x"f320";
    tmp(23299) := x"f300";
    tmp(23300) := x"eb00";
    tmp(23301) := x"f300";
    tmp(23302) := x"fb00";
    tmp(23303) := x"f320";
    tmp(23304) := x"f320";
    tmp(23305) := x"f340";
    tmp(23306) := x"f340";
    tmp(23307) := x"eb00";
    tmp(23308) := x"eae0";
    tmp(23309) := x"e2e0";
    tmp(23310) := x"dac0";
    tmp(23311) := x"c240";
    tmp(23312) := x"c260";
    tmp(23313) := x"e2e0";
    tmp(23314) := x"eb20";
    tmp(23315) := x"eb20";
    tmp(23316) := x"eb40";
    tmp(23317) := x"f360";
    tmp(23318) := x"f360";
    tmp(23319) := x"f380";
    tmp(23320) := x"fb80";
    tmp(23321) := x"f380";
    tmp(23322) := x"f380";
    tmp(23323) := x"fb80";
    tmp(23324) := x"eb40";
    tmp(23325) := x"eb40";
    tmp(23326) := x"eb40";
    tmp(23327) := x"eb40";
    tmp(23328) := x"fb60";
    tmp(23329) := x"fb80";
    tmp(23330) := x"fbe0";
    tmp(23331) := x"fbe0";
    tmp(23332) := x"fbc0";
    tmp(23333) := x"fbc0";
    tmp(23334) := x"fba0";
    tmp(23335) := x"fba0";
    tmp(23336) := x"fbc0";
    tmp(23337) := x"fbc0";
    tmp(23338) := x"fbc0";
    tmp(23339) := x"fba0";
    tmp(23340) := x"fb40";
    tmp(23341) := x"e2c0";
    tmp(23342) := x"e2a0";
    tmp(23343) := x"eaa0";
    tmp(23344) := x"eac0";
    tmp(23345) := x"f2e0";
    tmp(23346) := x"f300";
    tmp(23347) := x"fb60";
    tmp(23348) := x"fba0";
    tmp(23349) := x"fc40";
    tmp(23350) := x"fc40";
    tmp(23351) := x"fbe0";
    tmp(23352) := x"fb80";
    tmp(23353) := x"fb40";
    tmp(23354) := x"f300";
    tmp(23355) := x"f320";
    tmp(23356) := x"f320";
    tmp(23357) := x"f320";
    tmp(23358) := x"f320";
    tmp(23359) := x"f320";
    tmp(23360) := x"fb20";
    tmp(23361) := x"fb60";
    tmp(23362) := x"fba0";
    tmp(23363) := x"fba0";
    tmp(23364) := x"fb80";
    tmp(23365) := x"f300";
    tmp(23366) := x"eae0";
    tmp(23367) := x"f300";
    tmp(23368) := x"e2c0";
    tmp(23369) := x"dac0";
    tmp(23370) := x"f320";
    tmp(23371) := x"fb20";
    tmp(23372) := x"eae0";
    tmp(23373) := x"c240";
    tmp(23374) := x"b220";
    tmp(23375) := x"ba60";
    tmp(23376) := x"b240";
    tmp(23377) := x"99e0";
    tmp(23378) := x"91a0";
    tmp(23379) := x"99c0";
    tmp(23380) := x"99c0";
    tmp(23381) := x"99c0";
    tmp(23382) := x"a1c0";
    tmp(23383) := x"99c0";
    tmp(23384) := x"99c0";
    tmp(23385) := x"99e0";
    tmp(23386) := x"a200";
    tmp(23387) := x"9a00";
    tmp(23388) := x"b240";
    tmp(23389) := x"a220";
    tmp(23390) := x"9a40";
    tmp(23391) := x"69e0";
    tmp(23392) := x"2920";
    tmp(23393) := x"10e0";
    tmp(23394) := x"08c0";
    tmp(23395) := x"08c1";
    tmp(23396) := x"08c1";
    tmp(23397) := x"08c1";
    tmp(23398) := x"08a1";
    tmp(23399) := x"08c2";
    tmp(23400) := x"08c1";
    tmp(23401) := x"08e1";
    tmp(23402) := x"0902";
    tmp(23403) := x"0903";
    tmp(23404) := x"08e3";
    tmp(23405) := x"08c2";
    tmp(23406) := x"08e3";
    tmp(23407) := x"0924";
    tmp(23408) := x"0945";
    tmp(23409) := x"0965";
    tmp(23410) := x"0986";
    tmp(23411) := x"09a7";
    tmp(23412) := x"11e7";
    tmp(23413) := x"1aaa";
    tmp(23414) := x"1b2d";
    tmp(23415) := x"1b0c";
    tmp(23416) := x"33ae";
    tmp(23417) := x"8592";
    tmp(23418) := x"b5cf";
    tmp(23419) := x"b56d";
    tmp(23420) := x"b52d";
    tmp(23421) := x"b50c";
    tmp(23422) := x"b50c";
    tmp(23423) := x"aceb";
    tmp(23424) := x"9c6a";
    tmp(23425) := x"8be8";
    tmp(23426) := x"7ba8";
    tmp(23427) := x"6b46";
    tmp(23428) := x"6305";
    tmp(23429) := x"52a5";
    tmp(23430) := x"4264";
    tmp(23431) := x"3a43";
    tmp(23432) := x"31e2";
    tmp(23433) := x"31a2";
    tmp(23434) := x"31e2";
    tmp(23435) := x"4243";
    tmp(23436) := x"5ac4";
    tmp(23437) := x"6b45";
    tmp(23438) := x"83c7";
    tmp(23439) := x"a469";
    tmp(23440) := x"c52b";
    tmp(23441) := x"ddce";
    tmp(23442) := x"fed1";
    tmp(23443) := x"ff94";
    tmp(23444) := x"fff7";
    tmp(23445) := x"fffc";
    tmp(23446) := x"fffd";
    tmp(23447) := x"ffff";
    tmp(23448) := x"ffff";
    tmp(23449) := x"ffff";
    tmp(23450) := x"ffff";
    tmp(23451) := x"ffff";
    tmp(23452) := x"fffe";
    tmp(23453) := x"fffb";
    tmp(23454) := x"ff96";
    tmp(23455) := x"f691";
    tmp(23456) := x"ddee";
    tmp(23457) := x"c52d";
    tmp(23458) := x"93ea";
    tmp(23459) := x"7349";
    tmp(23460) := x"6b29";
    tmp(23461) := x"734b";
    tmp(23462) := x"7bac";
    tmp(23463) := x"940f";
    tmp(23464) := x"944f";
    tmp(23465) := x"9c71";
    tmp(23466) := x"9c72";
    tmp(23467) := x"ac92";
    tmp(23468) := x"bcf3";
    tmp(23469) := x"bcf4";
    tmp(23470) := x"bd15";
    tmp(23471) := x"bcf6";
    tmp(23472) := x"bd15";
    tmp(23473) := x"b4d4";
    tmp(23474) := x"ac95";
    tmp(23475) := x"a453";
    tmp(23476) := x"9c32";
    tmp(23477) := x"f800";
    tmp(23478) := x"f800";
    tmp(23479) := x"f800";
    tmp(23480) := x"f800";
    tmp(23481) := x"f800";
    tmp(23482) := x"f800";
    tmp(23483) := x"f800";
    tmp(23484) := x"f800";
    tmp(23485) := x"f800";
    tmp(23486) := x"f800";
    tmp(23487) := x"f800";
    tmp(23488) := x"f800";
    tmp(23489) := x"f800";
    tmp(23490) := x"f800";
    tmp(23491) := x"f800";
    tmp(23492) := x"f800";
    tmp(23493) := x"f800";
    tmp(23494) := x"f800";
    tmp(23495) := x"f800";
    tmp(23496) := x"f800";
    tmp(23497) := x"f800";
    tmp(23498) := x"f800";
    tmp(23499) := x"f800";
    tmp(23500) := x"f800";
    tmp(23501) := x"f800";
    tmp(23502) := x"f800";
    tmp(23503) := x"f800";
    tmp(23504) := x"f800";
    tmp(23505) := x"f800";
    tmp(23506) := x"f800";
    tmp(23507) := x"f800";
    tmp(23508) := x"f800";
    tmp(23509) := x"f800";
    tmp(23510) := x"f800";
    tmp(23511) := x"f800";
    tmp(23512) := x"f800";
    tmp(23513) := x"f800";
    tmp(23514) := x"f800";
    tmp(23515) := x"f800";
    tmp(23516) := x"f800";
    tmp(23517) := x"0840";
    tmp(23518) := x"0840";
    tmp(23519) := x"0840";
    tmp(23520) := x"1040";
    tmp(23521) := x"eb20";
    tmp(23522) := x"db00";
    tmp(23523) := x"eb40";
    tmp(23524) := x"f340";
    tmp(23525) := x"fb40";
    tmp(23526) := x"fb40";
    tmp(23527) := x"fb60";
    tmp(23528) := x"fb20";
    tmp(23529) := x"fb20";
    tmp(23530) := x"fb20";
    tmp(23531) := x"fb20";
    tmp(23532) := x"f2e0";
    tmp(23533) := x"fb20";
    tmp(23534) := x"fb40";
    tmp(23535) := x"fb20";
    tmp(23536) := x"fb40";
    tmp(23537) := x"fb40";
    tmp(23538) := x"fb20";
    tmp(23539) := x"f300";
    tmp(23540) := x"eae0";
    tmp(23541) := x"eae0";
    tmp(23542) := x"fb00";
    tmp(23543) := x"fb20";
    tmp(23544) := x"fb20";
    tmp(23545) := x"f340";
    tmp(23546) := x"fb40";
    tmp(23547) := x"eb00";
    tmp(23548) := x"f300";
    tmp(23549) := x"dac0";
    tmp(23550) := x"ca80";
    tmp(23551) := x"ca80";
    tmp(23552) := x"dac0";
    tmp(23553) := x"dae0";
    tmp(23554) := x"e300";
    tmp(23555) := x"eb20";
    tmp(23556) := x"eb40";
    tmp(23557) := x"eb40";
    tmp(23558) := x"eb40";
    tmp(23559) := x"fb80";
    tmp(23560) := x"fba0";
    tmp(23561) := x"fba0";
    tmp(23562) := x"fba0";
    tmp(23563) := x"f380";
    tmp(23564) := x"fb60";
    tmp(23565) := x"e320";
    tmp(23566) := x"e300";
    tmp(23567) := x"f340";
    tmp(23568) := x"f360";
    tmp(23569) := x"fb80";
    tmp(23570) := x"fbc0";
    tmp(23571) := x"fc00";
    tmp(23572) := x"fc00";
    tmp(23573) := x"fbc0";
    tmp(23574) := x"fb80";
    tmp(23575) := x"fb80";
    tmp(23576) := x"fba0";
    tmp(23577) := x"fba0";
    tmp(23578) := x"fb80";
    tmp(23579) := x"fba0";
    tmp(23580) := x"f320";
    tmp(23581) := x"fb00";
    tmp(23582) := x"eae0";
    tmp(23583) := x"eae0";
    tmp(23584) := x"e2a0";
    tmp(23585) := x"e280";
    tmp(23586) := x"fb20";
    tmp(23587) := x"f320";
    tmp(23588) := x"fb60";
    tmp(23589) := x"fbc0";
    tmp(23590) := x"fba0";
    tmp(23591) := x"fba0";
    tmp(23592) := x"fb60";
    tmp(23593) := x"fb60";
    tmp(23594) := x"fb40";
    tmp(23595) := x"fb20";
    tmp(23596) := x"fb40";
    tmp(23597) := x"fb40";
    tmp(23598) := x"fb60";
    tmp(23599) := x"fb60";
    tmp(23600) := x"fb40";
    tmp(23601) := x"fb80";
    tmp(23602) := x"fbc0";
    tmp(23603) := x"fbc0";
    tmp(23604) := x"fb80";
    tmp(23605) := x"fb60";
    tmp(23606) := x"fb40";
    tmp(23607) := x"f320";
    tmp(23608) := x"f300";
    tmp(23609) := x"eb20";
    tmp(23610) := x"fb40";
    tmp(23611) := x"fb20";
    tmp(23612) := x"f2e0";
    tmp(23613) := x"da80";
    tmp(23614) := x"c240";
    tmp(23615) := x"aa00";
    tmp(23616) := x"b200";
    tmp(23617) := x"a1e0";
    tmp(23618) := x"aa00";
    tmp(23619) := x"b200";
    tmp(23620) := x"aa00";
    tmp(23621) := x"a1e0";
    tmp(23622) := x"99c0";
    tmp(23623) := x"99e0";
    tmp(23624) := x"91e0";
    tmp(23625) := x"9a00";
    tmp(23626) := x"91c0";
    tmp(23627) := x"aa40";
    tmp(23628) := x"aa60";
    tmp(23629) := x"8a20";
    tmp(23630) := x"49a0";
    tmp(23631) := x"2120";
    tmp(23632) := x"10e0";
    tmp(23633) := x"08e0";
    tmp(23634) := x"0901";
    tmp(23635) := x"0901";
    tmp(23636) := x"08e2";
    tmp(23637) := x"08e2";
    tmp(23638) := x"08e2";
    tmp(23639) := x"08c2";
    tmp(23640) := x"08e2";
    tmp(23641) := x"0902";
    tmp(23642) := x"00c2";
    tmp(23643) := x"08c2";
    tmp(23644) := x"0903";
    tmp(23645) := x"08e3";
    tmp(23646) := x"0904";
    tmp(23647) := x"0945";
    tmp(23648) := x"09a6";
    tmp(23649) := x"09e8";
    tmp(23650) := x"126a";
    tmp(23651) := x"09c8";
    tmp(23652) := x"1229";
    tmp(23653) := x"122a";
    tmp(23654) := x"1a8b";
    tmp(23655) := x"3b4d";
    tmp(23656) := x"8d11";
    tmp(23657) := x"b5d0";
    tmp(23658) := x"bdae";
    tmp(23659) := x"bd6d";
    tmp(23660) := x"c56d";
    tmp(23661) := x"c54d";
    tmp(23662) := x"bd2c";
    tmp(23663) := x"bd2c";
    tmp(23664) := x"aceb";
    tmp(23665) := x"a48a";
    tmp(23666) := x"8be9";
    tmp(23667) := x"83a8";
    tmp(23668) := x"6b46";
    tmp(23669) := x"6326";
    tmp(23670) := x"5ac5";
    tmp(23671) := x"4a84";
    tmp(23672) := x"4243";
    tmp(23673) := x"3202";
    tmp(23674) := x"31c2";
    tmp(23675) := x"3a02";
    tmp(23676) := x"4a63";
    tmp(23677) := x"5ac4";
    tmp(23678) := x"7366";
    tmp(23679) := x"8be7";
    tmp(23680) := x"a48a";
    tmp(23681) := x"c56c";
    tmp(23682) := x"e60f";
    tmp(23683) := x"fe92";
    tmp(23684) := x"ffd5";
    tmp(23685) := x"fff7";
    tmp(23686) := x"fffd";
    tmp(23687) := x"ffff";
    tmp(23688) := x"ffff";
    tmp(23689) := x"ffff";
    tmp(23690) := x"ffff";
    tmp(23691) := x"ffff";
    tmp(23692) := x"ffff";
    tmp(23693) := x"fffc";
    tmp(23694) := x"fff8";
    tmp(23695) := x"fed2";
    tmp(23696) := x"edef";
    tmp(23697) := x"c52d";
    tmp(23698) := x"940a";
    tmp(23699) := x"7b69";
    tmp(23700) := x"734a";
    tmp(23701) := x"7b6c";
    tmp(23702) := x"83cd";
    tmp(23703) := x"8c0f";
    tmp(23704) := x"9c51";
    tmp(23705) := x"a492";
    tmp(23706) := x"acd3";
    tmp(23707) := x"acd3";
    tmp(23708) := x"acd3";
    tmp(23709) := x"bcf5";
    tmp(23710) := x"bd16";
    tmp(23711) := x"bcf6";
    tmp(23712) := x"c4f5";
    tmp(23713) := x"b4b4";
    tmp(23714) := x"ac94";
    tmp(23715) := x"ac74";
    tmp(23716) := x"9c53";
    tmp(23717) := x"f800";
    tmp(23718) := x"f800";
    tmp(23719) := x"f800";
    tmp(23720) := x"f800";
    tmp(23721) := x"f800";
    tmp(23722) := x"f800";
    tmp(23723) := x"f800";
    tmp(23724) := x"f800";
    tmp(23725) := x"f800";
    tmp(23726) := x"f800";
    tmp(23727) := x"f800";
    tmp(23728) := x"f800";
    tmp(23729) := x"f800";
    tmp(23730) := x"f800";
    tmp(23731) := x"f800";
    tmp(23732) := x"f800";
    tmp(23733) := x"f800";
    tmp(23734) := x"f800";
    tmp(23735) := x"f800";
    tmp(23736) := x"f800";
    tmp(23737) := x"f800";
    tmp(23738) := x"f800";
    tmp(23739) := x"f800";
    tmp(23740) := x"f800";
    tmp(23741) := x"f800";
    tmp(23742) := x"f800";
    tmp(23743) := x"f800";
    tmp(23744) := x"f800";
    tmp(23745) := x"f800";
    tmp(23746) := x"f800";
    tmp(23747) := x"f800";
    tmp(23748) := x"f800";
    tmp(23749) := x"f800";
    tmp(23750) := x"f800";
    tmp(23751) := x"f800";
    tmp(23752) := x"f800";
    tmp(23753) := x"f800";
    tmp(23754) := x"f800";
    tmp(23755) := x"f800";
    tmp(23756) := x"f800";
    tmp(23757) := x"0840";
    tmp(23758) := x"0840";
    tmp(23759) := x"0840";
    tmp(23760) := x"1040";
    tmp(23761) := x"dae0";
    tmp(23762) := x"dae0";
    tmp(23763) := x"eb20";
    tmp(23764) := x"eb00";
    tmp(23765) := x"f340";
    tmp(23766) := x"fb60";
    tmp(23767) := x"fb60";
    tmp(23768) := x"fb40";
    tmp(23769) := x"fb60";
    tmp(23770) := x"f320";
    tmp(23771) := x"f300";
    tmp(23772) := x"f300";
    tmp(23773) := x"f300";
    tmp(23774) := x"eae0";
    tmp(23775) := x"f320";
    tmp(23776) := x"f300";
    tmp(23777) := x"f300";
    tmp(23778) := x"f300";
    tmp(23779) := x"f300";
    tmp(23780) := x"f300";
    tmp(23781) := x"eae0";
    tmp(23782) := x"eae0";
    tmp(23783) := x"eb00";
    tmp(23784) := x"eb00";
    tmp(23785) := x"eb00";
    tmp(23786) := x"eb20";
    tmp(23787) := x"f320";
    tmp(23788) := x"e2e0";
    tmp(23789) := x"dac0";
    tmp(23790) := x"e2c0";
    tmp(23791) := x"d2a0";
    tmp(23792) := x"caa0";
    tmp(23793) := x"cac0";
    tmp(23794) := x"d2e0";
    tmp(23795) := x"db00";
    tmp(23796) := x"db20";
    tmp(23797) := x"db20";
    tmp(23798) := x"eb40";
    tmp(23799) := x"eb40";
    tmp(23800) := x"f360";
    tmp(23801) := x"fb80";
    tmp(23802) := x"fb80";
    tmp(23803) := x"fba0";
    tmp(23804) := x"fb60";
    tmp(23805) := x"eb40";
    tmp(23806) := x"e320";
    tmp(23807) := x"e300";
    tmp(23808) := x"fb60";
    tmp(23809) := x"fb80";
    tmp(23810) := x"fba0";
    tmp(23811) := x"fbc0";
    tmp(23812) := x"fbe0";
    tmp(23813) := x"fbc0";
    tmp(23814) := x"fba0";
    tmp(23815) := x"fba0";
    tmp(23816) := x"fbc0";
    tmp(23817) := x"fba0";
    tmp(23818) := x"fba0";
    tmp(23819) := x"fb40";
    tmp(23820) := x"f2e0";
    tmp(23821) := x"fb00";
    tmp(23822) := x"fb20";
    tmp(23823) := x"f2e0";
    tmp(23824) := x"eae0";
    tmp(23825) := x"eae0";
    tmp(23826) := x"eac0";
    tmp(23827) := x"f300";
    tmp(23828) := x"fb60";
    tmp(23829) := x"fba0";
    tmp(23830) := x"fba0";
    tmp(23831) := x"fb80";
    tmp(23832) := x"fbe0";
    tmp(23833) := x"fba0";
    tmp(23834) := x"fb40";
    tmp(23835) := x"fb20";
    tmp(23836) := x"fb80";
    tmp(23837) := x"fb80";
    tmp(23838) := x"fb80";
    tmp(23839) := x"fba0";
    tmp(23840) := x"fba0";
    tmp(23841) := x"fbc0";
    tmp(23842) := x"fbe0";
    tmp(23843) := x"fbc0";
    tmp(23844) := x"fb80";
    tmp(23845) := x"fb40";
    tmp(23846) := x"fb40";
    tmp(23847) := x"fb40";
    tmp(23848) := x"fb00";
    tmp(23849) := x"fb60";
    tmp(23850) := x"fb40";
    tmp(23851) := x"fb20";
    tmp(23852) := x"fb20";
    tmp(23853) := x"e2a0";
    tmp(23854) := x"ca60";
    tmp(23855) := x"b200";
    tmp(23856) := x"a9c0";
    tmp(23857) := x"a9e0";
    tmp(23858) := x"a9e0";
    tmp(23859) := x"b1e0";
    tmp(23860) := x"b200";
    tmp(23861) := x"a200";
    tmp(23862) := x"9a00";
    tmp(23863) := x"9a20";
    tmp(23864) := x"9a20";
    tmp(23865) := x"9a00";
    tmp(23866) := x"ba80";
    tmp(23867) := x"a260";
    tmp(23868) := x"61c0";
    tmp(23869) := x"3940";
    tmp(23870) := x"1920";
    tmp(23871) := x"08e0";
    tmp(23872) := x"08e1";
    tmp(23873) := x"08e1";
    tmp(23874) := x"08c1";
    tmp(23875) := x"08e1";
    tmp(23876) := x"08e1";
    tmp(23877) := x"0901";
    tmp(23878) := x"0902";
    tmp(23879) := x"0922";
    tmp(23880) := x"08e2";
    tmp(23881) := x"08e2";
    tmp(23882) := x"0922";
    tmp(23883) := x"0903";
    tmp(23884) := x"08e3";
    tmp(23885) := x"08e3";
    tmp(23886) := x"0945";
    tmp(23887) := x"0986";
    tmp(23888) := x"09a7";
    tmp(23889) := x"126a";
    tmp(23890) := x"1b4e";
    tmp(23891) := x"128c";
    tmp(23892) := x"1aac";
    tmp(23893) := x"22aa";
    tmp(23894) := x"3288";
    tmp(23895) := x"7c4c";
    tmp(23896) := x"94ad";
    tmp(23897) := x"a52d";
    tmp(23898) := x"b54d";
    tmp(23899) := x"c58d";
    tmp(23900) := x"c58d";
    tmp(23901) := x"cdad";
    tmp(23902) := x"c58d";
    tmp(23903) := x"c58d";
    tmp(23904) := x"c56d";
    tmp(23905) := x"b4eb";
    tmp(23906) := x"accb";
    tmp(23907) := x"9c4a";
    tmp(23908) := x"83a8";
    tmp(23909) := x"7387";
    tmp(23910) := x"6b26";
    tmp(23911) := x"5ae5";
    tmp(23912) := x"52a4";
    tmp(23913) := x"4263";
    tmp(23914) := x"3a22";
    tmp(23915) := x"31e2";
    tmp(23916) := x"4223";
    tmp(23917) := x"5284";
    tmp(23918) := x"6305";
    tmp(23919) := x"7b86";
    tmp(23920) := x"8c08";
    tmp(23921) := x"acea";
    tmp(23922) := x"cdac";
    tmp(23923) := x"ee90";
    tmp(23924) := x"ff12";
    tmp(23925) := x"ffd7";
    tmp(23926) := x"fff9";
    tmp(23927) := x"fffd";
    tmp(23928) := x"ffff";
    tmp(23929) := x"ffff";
    tmp(23930) := x"ffff";
    tmp(23931) := x"ffff";
    tmp(23932) := x"ffff";
    tmp(23933) := x"fffe";
    tmp(23934) := x"ffda";
    tmp(23935) := x"fef4";
    tmp(23936) := x"ee51";
    tmp(23937) := x"c52d";
    tmp(23938) := x"9c2b";
    tmp(23939) := x"7b4a";
    tmp(23940) := x"7b6b";
    tmp(23941) := x"8bce";
    tmp(23942) := x"93cf";
    tmp(23943) := x"940f";
    tmp(23944) := x"9c91";
    tmp(23945) := x"acd3";
    tmp(23946) := x"acd2";
    tmp(23947) := x"b4d3";
    tmp(23948) := x"b4d5";
    tmp(23949) := x"bcf5";
    tmp(23950) := x"bcf5";
    tmp(23951) := x"bd16";
    tmp(23952) := x"bcf5";
    tmp(23953) := x"b4b3";
    tmp(23954) := x"b4d5";
    tmp(23955) := x"a473";
    tmp(23956) := x"a473";
    tmp(23957) := x"f800";
    tmp(23958) := x"f800";
    tmp(23959) := x"f800";
    tmp(23960) := x"f800";
    tmp(23961) := x"f800";
    tmp(23962) := x"f800";
    tmp(23963) := x"f800";
    tmp(23964) := x"f800";
    tmp(23965) := x"f800";
    tmp(23966) := x"f800";
    tmp(23967) := x"f800";
    tmp(23968) := x"f800";
    tmp(23969) := x"f800";
    tmp(23970) := x"f800";
    tmp(23971) := x"f800";
    tmp(23972) := x"f800";
    tmp(23973) := x"f800";
    tmp(23974) := x"f800";
    tmp(23975) := x"f800";
    tmp(23976) := x"f800";
    tmp(23977) := x"f800";
    tmp(23978) := x"f800";
    tmp(23979) := x"f800";
    tmp(23980) := x"f800";
    tmp(23981) := x"f800";
    tmp(23982) := x"f800";
    tmp(23983) := x"f800";
    tmp(23984) := x"f800";
    tmp(23985) := x"f800";
    tmp(23986) := x"f800";
    tmp(23987) := x"f800";
    tmp(23988) := x"f800";
    tmp(23989) := x"f800";
    tmp(23990) := x"f800";
    tmp(23991) := x"f800";
    tmp(23992) := x"f800";
    tmp(23993) := x"f800";
    tmp(23994) := x"f800";
    tmp(23995) := x"f800";
    tmp(23996) := x"f800";
    tmp(23997) := x"0840";
    tmp(23998) := x"0840";
    tmp(23999) := x"0840";
    tmp(24000) := x"1040";
    tmp(24001) := x"e2e0";
    tmp(24002) := x"d2c0";
    tmp(24003) := x"db00";
    tmp(24004) := x"eb20";
    tmp(24005) := x"eb40";
    tmp(24006) := x"eb40";
    tmp(24007) := x"fb60";
    tmp(24008) := x"f340";
    tmp(24009) := x"f320";
    tmp(24010) := x"fb20";
    tmp(24011) := x"fb40";
    tmp(24012) := x"f300";
    tmp(24013) := x"f320";
    tmp(24014) := x"f300";
    tmp(24015) := x"f320";
    tmp(24016) := x"f300";
    tmp(24017) := x"f300";
    tmp(24018) := x"eae0";
    tmp(24019) := x"eb00";
    tmp(24020) := x"eae0";
    tmp(24021) := x"eb00";
    tmp(24022) := x"eae0";
    tmp(24023) := x"e2a0";
    tmp(24024) := x"e2c0";
    tmp(24025) := x"eae0";
    tmp(24026) := x"eb00";
    tmp(24027) := x"eb00";
    tmp(24028) := x"eb00";
    tmp(24029) := x"e2e0";
    tmp(24030) := x"dac0";
    tmp(24031) := x"d2a0";
    tmp(24032) := x"d2a0";
    tmp(24033) := x"ca80";
    tmp(24034) := x"cac0";
    tmp(24035) := x"e320";
    tmp(24036) := x"db20";
    tmp(24037) := x"db20";
    tmp(24038) := x"db20";
    tmp(24039) := x"e340";
    tmp(24040) := x"eb40";
    tmp(24041) := x"eb40";
    tmp(24042) := x"eb40";
    tmp(24043) := x"fba0";
    tmp(24044) := x"eb60";
    tmp(24045) := x"e320";
    tmp(24046) := x"dae0";
    tmp(24047) := x"fb60";
    tmp(24048) := x"f340";
    tmp(24049) := x"eb40";
    tmp(24050) := x"fba0";
    tmp(24051) := x"fb80";
    tmp(24052) := x"fba0";
    tmp(24053) := x"fba0";
    tmp(24054) := x"fba0";
    tmp(24055) := x"fba0";
    tmp(24056) := x"fba0";
    tmp(24057) := x"fba0";
    tmp(24058) := x"fba0";
    tmp(24059) := x"eb00";
    tmp(24060) := x"fb40";
    tmp(24061) := x"f300";
    tmp(24062) := x"fb80";
    tmp(24063) := x"fb80";
    tmp(24064) := x"f340";
    tmp(24065) := x"eb00";
    tmp(24066) := x"f2e0";
    tmp(24067) := x"f320";
    tmp(24068) := x"fb40";
    tmp(24069) := x"fb60";
    tmp(24070) := x"fb80";
    tmp(24071) := x"fc00";
    tmp(24072) := x"fc00";
    tmp(24073) := x"fba0";
    tmp(24074) := x"fb40";
    tmp(24075) := x"fb60";
    tmp(24076) := x"fb80";
    tmp(24077) := x"fba0";
    tmp(24078) := x"fb80";
    tmp(24079) := x"fbc0";
    tmp(24080) := x"fc20";
    tmp(24081) := x"fc40";
    tmp(24082) := x"fc20";
    tmp(24083) := x"fbe0";
    tmp(24084) := x"fb60";
    tmp(24085) := x"fb60";
    tmp(24086) := x"fb60";
    tmp(24087) := x"fb60";
    tmp(24088) := x"fb20";
    tmp(24089) := x"fb60";
    tmp(24090) := x"fb60";
    tmp(24091) := x"fb20";
    tmp(24092) := x"fb20";
    tmp(24093) := x"fb20";
    tmp(24094) := x"e2c0";
    tmp(24095) := x"c240";
    tmp(24096) := x"b220";
    tmp(24097) := x"a9e0";
    tmp(24098) := x"a1c0";
    tmp(24099) := x"aa00";
    tmp(24100) := x"9a00";
    tmp(24101) := x"9a40";
    tmp(24102) := x"bac0";
    tmp(24103) := x"a260";
    tmp(24104) := x"9220";
    tmp(24105) := x"9a40";
    tmp(24106) := x"9a20";
    tmp(24107) := x"5160";
    tmp(24108) := x"2100";
    tmp(24109) := x"10e0";
    tmp(24110) := x"08e0";
    tmp(24111) := x"0901";
    tmp(24112) := x"0901";
    tmp(24113) := x"0901";
    tmp(24114) := x"08e1";
    tmp(24115) := x"08e1";
    tmp(24116) := x"08c1";
    tmp(24117) := x"08a0";
    tmp(24118) := x"0901";
    tmp(24119) := x"0922";
    tmp(24120) := x"0902";
    tmp(24121) := x"0902";
    tmp(24122) := x"0943";
    tmp(24123) := x"0944";
    tmp(24124) := x"0965";
    tmp(24125) := x"0985";
    tmp(24126) := x"09a7";
    tmp(24127) := x"0986";
    tmp(24128) := x"11e8";
    tmp(24129) := x"1acd";
    tmp(24130) := x"1acd";
    tmp(24131) := x"22ed";
    tmp(24132) := x"2268";
    tmp(24133) := x"3245";
    tmp(24134) := x"5307";
    tmp(24135) := x"6b47";
    tmp(24136) := x"7bc9";
    tmp(24137) := x"946b";
    tmp(24138) := x"a4ec";
    tmp(24139) := x"b50d";
    tmp(24140) := x"bd2d";
    tmp(24141) := x"cd8d";
    tmp(24142) := x"cdce";
    tmp(24143) := x"cdae";
    tmp(24144) := x"cdce";
    tmp(24145) := x"c56d";
    tmp(24146) := x"bd4c";
    tmp(24147) := x"accb";
    tmp(24148) := x"946a";
    tmp(24149) := x"8c09";
    tmp(24150) := x"7b67";
    tmp(24151) := x"6b26";
    tmp(24152) := x"5ae5";
    tmp(24153) := x"52c4";
    tmp(24154) := x"4a64";
    tmp(24155) := x"4243";
    tmp(24156) := x"3a02";
    tmp(24157) := x"4243";
    tmp(24158) := x"52a4";
    tmp(24159) := x"6b45";
    tmp(24160) := x"7ba6";
    tmp(24161) := x"9448";
    tmp(24162) := x"bd0b";
    tmp(24163) := x"cdae";
    tmp(24164) := x"fef1";
    tmp(24165) := x"ff74";
    tmp(24166) := x"ffd8";
    tmp(24167) := x"fffa";
    tmp(24168) := x"fffe";
    tmp(24169) := x"ffff";
    tmp(24170) := x"ffff";
    tmp(24171) := x"ffff";
    tmp(24172) := x"ffff";
    tmp(24173) := x"fffe";
    tmp(24174) := x"fff9";
    tmp(24175) := x"ff55";
    tmp(24176) := x"feb2";
    tmp(24177) := x"cd6e";
    tmp(24178) := x"9c2c";
    tmp(24179) := x"836a";
    tmp(24180) := x"836c";
    tmp(24181) := x"8bce";
    tmp(24182) := x"940f";
    tmp(24183) := x"9c71";
    tmp(24184) := x"acd2";
    tmp(24185) := x"b4f3";
    tmp(24186) := x"bd55";
    tmp(24187) := x"bd36";
    tmp(24188) := x"b515";
    tmp(24189) := x"bd15";
    tmp(24190) := x"bcd5";
    tmp(24191) := x"c516";
    tmp(24192) := x"bcf5";
    tmp(24193) := x"b4d4";
    tmp(24194) := x"b4d4";
    tmp(24195) := x"ac94";
    tmp(24196) := x"acd4";
    tmp(24197) := x"f800";
    tmp(24198) := x"f800";
    tmp(24199) := x"f800";
    tmp(24200) := x"f800";
    tmp(24201) := x"f800";
    tmp(24202) := x"f800";
    tmp(24203) := x"f800";
    tmp(24204) := x"f800";
    tmp(24205) := x"f800";
    tmp(24206) := x"f800";
    tmp(24207) := x"f800";
    tmp(24208) := x"f800";
    tmp(24209) := x"f800";
    tmp(24210) := x"f800";
    tmp(24211) := x"f800";
    tmp(24212) := x"f800";
    tmp(24213) := x"f800";
    tmp(24214) := x"f800";
    tmp(24215) := x"f800";
    tmp(24216) := x"f800";
    tmp(24217) := x"f800";
    tmp(24218) := x"f800";
    tmp(24219) := x"f800";
    tmp(24220) := x"f800";
    tmp(24221) := x"f800";
    tmp(24222) := x"f800";
    tmp(24223) := x"f800";
    tmp(24224) := x"f800";
    tmp(24225) := x"f800";
    tmp(24226) := x"f800";
    tmp(24227) := x"f800";
    tmp(24228) := x"f800";
    tmp(24229) := x"f800";
    tmp(24230) := x"f800";
    tmp(24231) := x"f800";
    tmp(24232) := x"f800";
    tmp(24233) := x"f800";
    tmp(24234) := x"f800";
    tmp(24235) := x"f800";
    tmp(24236) := x"f800";
    tmp(24237) := x"0840";
    tmp(24238) := x"0840";
    tmp(24239) := x"0840";
    tmp(24240) := x"1040";
    tmp(24241) := x"dac0";
    tmp(24242) := x"caa0";
    tmp(24243) := x"cac0";
    tmp(24244) := x"dac0";
    tmp(24245) := x"e320";
    tmp(24246) := x"f340";
    tmp(24247) := x"eb20";
    tmp(24248) := x"eb00";
    tmp(24249) := x"fb20";
    tmp(24250) := x"fb00";
    tmp(24251) := x"f320";
    tmp(24252) := x"eb00";
    tmp(24253) := x"f320";
    tmp(24254) := x"eb00";
    tmp(24255) := x"eb00";
    tmp(24256) := x"eae0";
    tmp(24257) := x"e2c0";
    tmp(24258) := x"dac0";
    tmp(24259) := x"dac0";
    tmp(24260) := x"e2c0";
    tmp(24261) := x"e2c0";
    tmp(24262) := x"dac0";
    tmp(24263) := x"daa0";
    tmp(24264) := x"d2a0";
    tmp(24265) := x"dac0";
    tmp(24266) := x"e2c0";
    tmp(24267) := x"dac0";
    tmp(24268) := x"dac0";
    tmp(24269) := x"daa0";
    tmp(24270) := x"d2a0";
    tmp(24271) := x"d2c0";
    tmp(24272) := x"caa0";
    tmp(24273) := x"caa0";
    tmp(24274) := x"d2e0";
    tmp(24275) := x"d2e0";
    tmp(24276) := x"d300";
    tmp(24277) := x"d300";
    tmp(24278) := x"db00";
    tmp(24279) := x"e340";
    tmp(24280) := x"eb40";
    tmp(24281) := x"eb60";
    tmp(24282) := x"eb60";
    tmp(24283) := x"eb60";
    tmp(24284) := x"d2e0";
    tmp(24285) := x"db00";
    tmp(24286) := x"e340";
    tmp(24287) := x"db20";
    tmp(24288) := x"e300";
    tmp(24289) := x"eb40";
    tmp(24290) := x"f380";
    tmp(24291) := x"f360";
    tmp(24292) := x"f380";
    tmp(24293) := x"fb80";
    tmp(24294) := x"fbc0";
    tmp(24295) := x"fbe0";
    tmp(24296) := x"fbe0";
    tmp(24297) := x"fbc0";
    tmp(24298) := x"fba0";
    tmp(24299) := x"fb80";
    tmp(24300) := x"eb20";
    tmp(24301) := x"fb60";
    tmp(24302) := x"fb80";
    tmp(24303) := x"fb80";
    tmp(24304) := x"f360";
    tmp(24305) := x"dac0";
    tmp(24306) := x"dac0";
    tmp(24307) := x"e2e0";
    tmp(24308) := x"e2c0";
    tmp(24309) := x"fb40";
    tmp(24310) := x"fbc0";
    tmp(24311) := x"fbe0";
    tmp(24312) := x"fc00";
    tmp(24313) := x"fbc0";
    tmp(24314) := x"fb80";
    tmp(24315) := x"fba0";
    tmp(24316) := x"f340";
    tmp(24317) := x"fb60";
    tmp(24318) := x"fba0";
    tmp(24319) := x"fbe0";
    tmp(24320) := x"fc00";
    tmp(24321) := x"fc20";
    tmp(24322) := x"fc00";
    tmp(24323) := x"fbe0";
    tmp(24324) := x"fba0";
    tmp(24325) := x"fb80";
    tmp(24326) := x"fb80";
    tmp(24327) := x"fb40";
    tmp(24328) := x"fb60";
    tmp(24329) := x"fb00";
    tmp(24330) := x"f2e0";
    tmp(24331) := x"fb40";
    tmp(24332) := x"fb40";
    tmp(24333) := x"f340";
    tmp(24334) := x"f340";
    tmp(24335) := x"c240";
    tmp(24336) := x"99c0";
    tmp(24337) := x"91c0";
    tmp(24338) := x"91e0";
    tmp(24339) := x"8a00";
    tmp(24340) := x"9240";
    tmp(24341) := x"a2a0";
    tmp(24342) := x"9a80";
    tmp(24343) := x"8220";
    tmp(24344) := x"79e0";
    tmp(24345) := x"8200";
    tmp(24346) := x"7a00";
    tmp(24347) := x"49a0";
    tmp(24348) := x"10e0";
    tmp(24349) := x"08c0";
    tmp(24350) := x"08c1";
    tmp(24351) := x"08e1";
    tmp(24352) := x"08e1";
    tmp(24353) := x"08c0";
    tmp(24354) := x"08c0";
    tmp(24355) := x"08e1";
    tmp(24356) := x"0901";
    tmp(24357) := x"08e1";
    tmp(24358) := x"0942";
    tmp(24359) := x"0943";
    tmp(24360) := x"0922";
    tmp(24361) := x"0964";
    tmp(24362) := x"0986";
    tmp(24363) := x"0966";
    tmp(24364) := x"09a7";
    tmp(24365) := x"09a7";
    tmp(24366) := x"11e8";
    tmp(24367) := x"1229";
    tmp(24368) := x"1a8b";
    tmp(24369) := x"230d";
    tmp(24370) := x"2acb";
    tmp(24371) := x"21e6";
    tmp(24372) := x"21a4";
    tmp(24373) := x"3203";
    tmp(24374) := x"4244";
    tmp(24375) := x"52c5";
    tmp(24376) := x"5b27";
    tmp(24377) := x"6b68";
    tmp(24378) := x"83ea";
    tmp(24379) := x"9c8b";
    tmp(24380) := x"bd4d";
    tmp(24381) := x"c58d";
    tmp(24382) := x"cdad";
    tmp(24383) := x"d5ee";
    tmp(24384) := x"ddee";
    tmp(24385) := x"cdee";
    tmp(24386) := x"d5ee";
    tmp(24387) := x"c56d";
    tmp(24388) := x"aceb";
    tmp(24389) := x"9c6a";
    tmp(24390) := x"942a";
    tmp(24391) := x"7b88";
    tmp(24392) := x"7347";
    tmp(24393) := x"5b05";
    tmp(24394) := x"52c5";
    tmp(24395) := x"4a84";
    tmp(24396) := x"4243";
    tmp(24397) := x"3a43";
    tmp(24398) := x"4263";
    tmp(24399) := x"52c4";
    tmp(24400) := x"6b46";
    tmp(24401) := x"83c7";
    tmp(24402) := x"9c69";
    tmp(24403) := x"bd4d";
    tmp(24404) := x"e60e";
    tmp(24405) := x"f691";
    tmp(24406) := x"ffb5";
    tmp(24407) := x"fff8";
    tmp(24408) := x"fffb";
    tmp(24409) := x"fffd";
    tmp(24410) := x"ffff";
    tmp(24411) := x"ffff";
    tmp(24412) := x"ffff";
    tmp(24413) := x"fffe";
    tmp(24414) := x"fffa";
    tmp(24415) := x"ff35";
    tmp(24416) := x"feb3";
    tmp(24417) := x"d58f";
    tmp(24418) := x"9c0c";
    tmp(24419) := x"8bcc";
    tmp(24420) := x"93ee";
    tmp(24421) := x"940f";
    tmp(24422) := x"9c70";
    tmp(24423) := x"a492";
    tmp(24424) := x"a4b2";
    tmp(24425) := x"acb3";
    tmp(24426) := x"b4f5";
    tmp(24427) := x"b4f4";
    tmp(24428) := x"b4f4";
    tmp(24429) := x"bcf5";
    tmp(24430) := x"bcf6";
    tmp(24431) := x"b4f5";
    tmp(24432) := x"bcf4";
    tmp(24433) := x"b4f5";
    tmp(24434) := x"bcf6";
    tmp(24435) := x"b4d5";
    tmp(24436) := x"ac74";
    tmp(24437) := x"f800";
    tmp(24438) := x"f800";
    tmp(24439) := x"f800";
    tmp(24440) := x"f800";
    tmp(24441) := x"f800";
    tmp(24442) := x"f800";
    tmp(24443) := x"f800";
    tmp(24444) := x"f800";
    tmp(24445) := x"f800";
    tmp(24446) := x"f800";
    tmp(24447) := x"f800";
    tmp(24448) := x"f800";
    tmp(24449) := x"f800";
    tmp(24450) := x"f800";
    tmp(24451) := x"f800";
    tmp(24452) := x"f800";
    tmp(24453) := x"f800";
    tmp(24454) := x"f800";
    tmp(24455) := x"f800";
    tmp(24456) := x"f800";
    tmp(24457) := x"f800";
    tmp(24458) := x"f800";
    tmp(24459) := x"f800";
    tmp(24460) := x"f800";
    tmp(24461) := x"f800";
    tmp(24462) := x"f800";
    tmp(24463) := x"f800";
    tmp(24464) := x"f800";
    tmp(24465) := x"f800";
    tmp(24466) := x"f800";
    tmp(24467) := x"f800";
    tmp(24468) := x"f800";
    tmp(24469) := x"f800";
    tmp(24470) := x"f800";
    tmp(24471) := x"f800";
    tmp(24472) := x"f800";
    tmp(24473) := x"f800";
    tmp(24474) := x"f800";
    tmp(24475) := x"f800";
    tmp(24476) := x"f800";
    tmp(24477) := x"0840";
    tmp(24478) := x"0840";
    tmp(24479) := x"0840";
    tmp(24480) := x"1040";
    tmp(24481) := x"caa0";
    tmp(24482) := x"c280";
    tmp(24483) := x"c280";
    tmp(24484) := x"cac0";
    tmp(24485) := x"d2c0";
    tmp(24486) := x"e300";
    tmp(24487) := x"dae0";
    tmp(24488) := x"e2e0";
    tmp(24489) := x"e2c0";
    tmp(24490) := x"eac0";
    tmp(24491) := x"eae0";
    tmp(24492) := x"eae0";
    tmp(24493) := x"f320";
    tmp(24494) := x"eb00";
    tmp(24495) := x"eb00";
    tmp(24496) := x"eb00";
    tmp(24497) := x"daa0";
    tmp(24498) := x"d2a0";
    tmp(24499) := x"ca80";
    tmp(24500) := x"d2a0";
    tmp(24501) := x"e2c0";
    tmp(24502) := x"d2a0";
    tmp(24503) := x"ca80";
    tmp(24504) := x"ca80";
    tmp(24505) := x"c260";
    tmp(24506) := x"c260";
    tmp(24507) := x"ca80";
    tmp(24508) := x"c280";
    tmp(24509) := x"ca80";
    tmp(24510) := x"c280";
    tmp(24511) := x"cac0";
    tmp(24512) := x"caa0";
    tmp(24513) := x"cac0";
    tmp(24514) := x"cac0";
    tmp(24515) := x"cac0";
    tmp(24516) := x"c2c0";
    tmp(24517) := x"cac0";
    tmp(24518) := x"d300";
    tmp(24519) := x"db20";
    tmp(24520) := x"db20";
    tmp(24521) := x"db20";
    tmp(24522) := x"d320";
    tmp(24523) := x"d320";
    tmp(24524) := x"cac0";
    tmp(24525) := x"b260";
    tmp(24526) := x"cb00";
    tmp(24527) := x"db20";
    tmp(24528) := x"d2e0";
    tmp(24529) := x"eb60";
    tmp(24530) := x"db20";
    tmp(24531) := x"eb40";
    tmp(24532) := x"eb60";
    tmp(24533) := x"f360";
    tmp(24534) := x"eb60";
    tmp(24535) := x"fbc0";
    tmp(24536) := x"fbe0";
    tmp(24537) := x"fbc0";
    tmp(24538) := x"fbc0";
    tmp(24539) := x"fbc0";
    tmp(24540) := x"fbc0";
    tmp(24541) := x"eb40";
    tmp(24542) := x"f320";
    tmp(24543) := x"fb60";
    tmp(24544) := x"eb40";
    tmp(24545) := x"e300";
    tmp(24546) := x"d2a0";
    tmp(24547) := x"c240";
    tmp(24548) := x"e2c0";
    tmp(24549) := x"fb60";
    tmp(24550) := x"fb80";
    tmp(24551) := x"fbc0";
    tmp(24552) := x"fbe0";
    tmp(24553) := x"fc00";
    tmp(24554) := x"fc20";
    tmp(24555) := x"fb80";
    tmp(24556) := x"fba0";
    tmp(24557) := x"fba0";
    tmp(24558) := x"fbc0";
    tmp(24559) := x"fc00";
    tmp(24560) := x"fbe0";
    tmp(24561) := x"fbc0";
    tmp(24562) := x"fbc0";
    tmp(24563) := x"fba0";
    tmp(24564) := x"fbc0";
    tmp(24565) := x"fbc0";
    tmp(24566) := x"fbe0";
    tmp(24567) := x"fbc0";
    tmp(24568) := x"fb60";
    tmp(24569) := x"fb40";
    tmp(24570) := x"f320";
    tmp(24571) := x"fb40";
    tmp(24572) := x"f320";
    tmp(24573) := x"fb60";
    tmp(24574) := x"eae0";
    tmp(24575) := x"b220";
    tmp(24576) := x"89a0";
    tmp(24577) := x"6980";
    tmp(24578) := x"6180";
    tmp(24579) := x"71e0";
    tmp(24580) := x"8240";
    tmp(24581) := x"7a40";
    tmp(24582) := x"61c0";
    tmp(24583) := x"5180";
    tmp(24584) := x"5180";
    tmp(24585) := x"6a00";
    tmp(24586) := x"51e0";
    tmp(24587) := x"2121";
    tmp(24588) := x"08e1";
    tmp(24589) := x"08a1";
    tmp(24590) := x"08c1";
    tmp(24591) := x"0901";
    tmp(24592) := x"08e1";
    tmp(24593) := x"08e1";
    tmp(24594) := x"08e1";
    tmp(24595) := x"0921";
    tmp(24596) := x"0942";
    tmp(24597) := x"0942";
    tmp(24598) := x"0902";
    tmp(24599) := x"0923";
    tmp(24600) := x"0903";
    tmp(24601) := x"0965";
    tmp(24602) := x"09a7";
    tmp(24603) := x"11e8";
    tmp(24604) := x"1209";
    tmp(24605) := x"1229";
    tmp(24606) := x"1aab";
    tmp(24607) := x"2b8e";
    tmp(24608) := x"442f";
    tmp(24609) := x"436b";
    tmp(24610) := x"3a47";
    tmp(24611) := x"29e5";
    tmp(24612) := x"29a4";
    tmp(24613) := x"2183";
    tmp(24614) := x"29c2";
    tmp(24615) := x"3a23";
    tmp(24616) := x"4a84";
    tmp(24617) := x"5b06";
    tmp(24618) := x"6b67";
    tmp(24619) := x"83c9";
    tmp(24620) := x"9c8a";
    tmp(24621) := x"b52c";
    tmp(24622) := x"c58c";
    tmp(24623) := x"d5cd";
    tmp(24624) := x"de0e";
    tmp(24625) := x"de2f";
    tmp(24626) := x"de10";
    tmp(24627) := x"cdae";
    tmp(24628) := x"bd6d";
    tmp(24629) := x"b4cc";
    tmp(24630) := x"a46b";
    tmp(24631) := x"9429";
    tmp(24632) := x"7ba8";
    tmp(24633) := x"7347";
    tmp(24634) := x"6326";
    tmp(24635) := x"52c5";
    tmp(24636) := x"4a84";
    tmp(24637) := x"4243";
    tmp(24638) := x"3a43";
    tmp(24639) := x"4a83";
    tmp(24640) := x"5ae4";
    tmp(24641) := x"6b46";
    tmp(24642) := x"83c7";
    tmp(24643) := x"a489";
    tmp(24644) := x"bd2c";
    tmp(24645) := x"e5ef";
    tmp(24646) := x"f6d1";
    tmp(24647) := x"ff95";
    tmp(24648) := x"fff9";
    tmp(24649) := x"fffd";
    tmp(24650) := x"fffe";
    tmp(24651) := x"ffff";
    tmp(24652) := x"ffff";
    tmp(24653) := x"ffff";
    tmp(24654) := x"fffc";
    tmp(24655) := x"ff97";
    tmp(24656) := x"fed4";
    tmp(24657) := x"ddb1";
    tmp(24658) := x"ac8e";
    tmp(24659) := x"93ed";
    tmp(24660) := x"93ce";
    tmp(24661) := x"9c50";
    tmp(24662) := x"a471";
    tmp(24663) := x"acd3";
    tmp(24664) := x"acd4";
    tmp(24665) := x"b4f5";
    tmp(24666) := x"b4d5";
    tmp(24667) := x"b515";
    tmp(24668) := x"bd35";
    tmp(24669) := x"bd16";
    tmp(24670) := x"c516";
    tmp(24671) := x"bd17";
    tmp(24672) := x"b4d5";
    tmp(24673) := x"bcf5";
    tmp(24674) := x"b494";
    tmp(24675) := x"ac94";
    tmp(24676) := x"b4b4";
    tmp(24677) := x"f800";
    tmp(24678) := x"f800";
    tmp(24679) := x"f800";
    tmp(24680) := x"f800";
    tmp(24681) := x"f800";
    tmp(24682) := x"f800";
    tmp(24683) := x"f800";
    tmp(24684) := x"f800";
    tmp(24685) := x"f800";
    tmp(24686) := x"f800";
    tmp(24687) := x"f800";
    tmp(24688) := x"f800";
    tmp(24689) := x"f800";
    tmp(24690) := x"f800";
    tmp(24691) := x"f800";
    tmp(24692) := x"f800";
    tmp(24693) := x"f800";
    tmp(24694) := x"f800";
    tmp(24695) := x"f800";
    tmp(24696) := x"f800";
    tmp(24697) := x"f800";
    tmp(24698) := x"f800";
    tmp(24699) := x"f800";
    tmp(24700) := x"f800";
    tmp(24701) := x"f800";
    tmp(24702) := x"f800";
    tmp(24703) := x"f800";
    tmp(24704) := x"f800";
    tmp(24705) := x"f800";
    tmp(24706) := x"f800";
    tmp(24707) := x"f800";
    tmp(24708) := x"f800";
    tmp(24709) := x"f800";
    tmp(24710) := x"f800";
    tmp(24711) := x"f800";
    tmp(24712) := x"f800";
    tmp(24713) := x"f800";
    tmp(24714) := x"f800";
    tmp(24715) := x"f800";
    tmp(24716) := x"f800";
    tmp(24717) := x"0840";
    tmp(24718) := x"0840";
    tmp(24719) := x"0840";
    tmp(24720) := x"1040";
    tmp(24721) := x"ba80";
    tmp(24722) := x"ba80";
    tmp(24723) := x"b280";
    tmp(24724) := x"ba80";
    tmp(24725) := x"cac0";
    tmp(24726) := x"d2c0";
    tmp(24727) := x"caa0";
    tmp(24728) := x"dac0";
    tmp(24729) := x"e2c0";
    tmp(24730) := x"e2c0";
    tmp(24731) := x"e2e0";
    tmp(24732) := x"e2e0";
    tmp(24733) := x"eb00";
    tmp(24734) := x"e2e0";
    tmp(24735) := x"eb00";
    tmp(24736) := x"dae0";
    tmp(24737) := x"ca80";
    tmp(24738) := x"d280";
    tmp(24739) := x"ca80";
    tmp(24740) := x"ca80";
    tmp(24741) := x"d280";
    tmp(24742) := x"ca80";
    tmp(24743) := x"caa0";
    tmp(24744) := x"c280";
    tmp(24745) := x"ba40";
    tmp(24746) := x"b240";
    tmp(24747) := x"b220";
    tmp(24748) := x"ba60";
    tmp(24749) := x"ba60";
    tmp(24750) := x"caa0";
    tmp(24751) := x"ba80";
    tmp(24752) := x"c2a0";
    tmp(24753) := x"b260";
    tmp(24754) := x"b280";
    tmp(24755) := x"b280";
    tmp(24756) := x"bac0";
    tmp(24757) := x"c2e0";
    tmp(24758) := x"cae0";
    tmp(24759) := x"c2c0";
    tmp(24760) := x"c2e0";
    tmp(24761) := x"c2e0";
    tmp(24762) := x"c2c0";
    tmp(24763) := x"c2e0";
    tmp(24764) := x"aa60";
    tmp(24765) := x"b2c0";
    tmp(24766) := x"bac0";
    tmp(24767) := x"c2c0";
    tmp(24768) := x"cae0";
    tmp(24769) := x"cb00";
    tmp(24770) := x"d340";
    tmp(24771) := x"db20";
    tmp(24772) := x"e340";
    tmp(24773) := x"eb60";
    tmp(24774) := x"f3c0";
    tmp(24775) := x"f3c0";
    tmp(24776) := x"eba0";
    tmp(24777) := x"fbe0";
    tmp(24778) := x"fc60";
    tmp(24779) := x"eba0";
    tmp(24780) := x"eb80";
    tmp(24781) := x"d300";
    tmp(24782) := x"dae0";
    tmp(24783) := x"e320";
    tmp(24784) := x"eb40";
    tmp(24785) := x"dae0";
    tmp(24786) := x"d2c0";
    tmp(24787) := x"d2a0";
    tmp(24788) := x"dac0";
    tmp(24789) := x"f320";
    tmp(24790) := x"fb40";
    tmp(24791) := x"fbc0";
    tmp(24792) := x"fbe0";
    tmp(24793) := x"fbe0";
    tmp(24794) := x"fba0";
    tmp(24795) := x"f3a0";
    tmp(24796) := x"f380";
    tmp(24797) := x"eb60";
    tmp(24798) := x"fc00";
    tmp(24799) := x"fb80";
    tmp(24800) := x"fba0";
    tmp(24801) := x"f380";
    tmp(24802) := x"fb80";
    tmp(24803) := x"fba0";
    tmp(24804) := x"fbc0";
    tmp(24805) := x"fc00";
    tmp(24806) := x"fbe0";
    tmp(24807) := x"fc00";
    tmp(24808) := x"fba0";
    tmp(24809) := x"eb00";
    tmp(24810) := x"fb60";
    tmp(24811) := x"f320";
    tmp(24812) := x"eb40";
    tmp(24813) := x"f340";
    tmp(24814) := x"e2e0";
    tmp(24815) := x"a200";
    tmp(24816) := x"5980";
    tmp(24817) := x"4140";
    tmp(24818) := x"4980";
    tmp(24819) := x"49a0";
    tmp(24820) := x"4980";
    tmp(24821) := x"3940";
    tmp(24822) := x"3940";
    tmp(24823) := x"3960";
    tmp(24824) := x"3980";
    tmp(24825) := x"2161";
    tmp(24826) := x"1122";
    tmp(24827) := x"08e2";
    tmp(24828) := x"0902";
    tmp(24829) := x"08c1";
    tmp(24830) := x"0901";
    tmp(24831) := x"0942";
    tmp(24832) := x"0901";
    tmp(24833) := x"0902";
    tmp(24834) := x"0922";
    tmp(24835) := x"0943";
    tmp(24836) := x"09a5";
    tmp(24837) := x"09c5";
    tmp(24838) := x"0984";
    tmp(24839) := x"11e6";
    tmp(24840) := x"09a6";
    tmp(24841) := x"0986";
    tmp(24842) := x"11e9";
    tmp(24843) := x"1209";
    tmp(24844) := x"1208";
    tmp(24845) := x"228a";
    tmp(24846) := x"43ce";
    tmp(24847) := x"6c4e";
    tmp(24848) := x"636a";
    tmp(24849) := x"5ae8";
    tmp(24850) := x"4aa8";
    tmp(24851) := x"3a67";
    tmp(24852) := x"3206";
    tmp(24853) := x"21a3";
    tmp(24854) := x"2162";
    tmp(24855) := x"2182";
    tmp(24856) := x"31e2";
    tmp(24857) := x"4244";
    tmp(24858) := x"52c5";
    tmp(24859) := x"6b47";
    tmp(24860) := x"83e8";
    tmp(24861) := x"9c89";
    tmp(24862) := x"b4ea";
    tmp(24863) := x"cdad";
    tmp(24864) := x"d5ee";
    tmp(24865) := x"de2f";
    tmp(24866) := x"e630";
    tmp(24867) := x"de30";
    tmp(24868) := x"d5ef";
    tmp(24869) := x"cd8e";
    tmp(24870) := x"b4ec";
    tmp(24871) := x"a48b";
    tmp(24872) := x"9409";
    tmp(24873) := x"83a8";
    tmp(24874) := x"7347";
    tmp(24875) := x"6306";
    tmp(24876) := x"5ac5";
    tmp(24877) := x"4a84";
    tmp(24878) := x"4264";
    tmp(24879) := x"4243";
    tmp(24880) := x"4a63";
    tmp(24881) := x"52c4";
    tmp(24882) := x"6b26";
    tmp(24883) := x"9408";
    tmp(24884) := x"9c6a";
    tmp(24885) := x"bd2d";
    tmp(24886) := x"ddef";
    tmp(24887) := x"f6d2";
    tmp(24888) := x"ff95";
    tmp(24889) := x"fff9";
    tmp(24890) := x"fffb";
    tmp(24891) := x"fffe";
    tmp(24892) := x"ffff";
    tmp(24893) := x"ffff";
    tmp(24894) := x"fffb";
    tmp(24895) := x"ff98";
    tmp(24896) := x"fef5";
    tmp(24897) := x"e612";
    tmp(24898) := x"ac8e";
    tmp(24899) := x"a44f";
    tmp(24900) := x"9c50";
    tmp(24901) := x"a471";
    tmp(24902) := x"b4d2";
    tmp(24903) := x"acb3";
    tmp(24904) := x"b4d4";
    tmp(24905) := x"b4f5";
    tmp(24906) := x"bd15";
    tmp(24907) := x"b515";
    tmp(24908) := x"b515";
    tmp(24909) := x"bcf6";
    tmp(24910) := x"bcf6";
    tmp(24911) := x"bcf6";
    tmp(24912) := x"bcf6";
    tmp(24913) := x"bcf6";
    tmp(24914) := x"bcd5";
    tmp(24915) := x"ac94";
    tmp(24916) := x"ac95";
    tmp(24917) := x"f800";
    tmp(24918) := x"f800";
    tmp(24919) := x"f800";
    tmp(24920) := x"f800";
    tmp(24921) := x"f800";
    tmp(24922) := x"f800";
    tmp(24923) := x"f800";
    tmp(24924) := x"f800";
    tmp(24925) := x"f800";
    tmp(24926) := x"f800";
    tmp(24927) := x"f800";
    tmp(24928) := x"f800";
    tmp(24929) := x"f800";
    tmp(24930) := x"f800";
    tmp(24931) := x"f800";
    tmp(24932) := x"f800";
    tmp(24933) := x"f800";
    tmp(24934) := x"f800";
    tmp(24935) := x"f800";
    tmp(24936) := x"f800";
    tmp(24937) := x"f800";
    tmp(24938) := x"f800";
    tmp(24939) := x"f800";
    tmp(24940) := x"f800";
    tmp(24941) := x"f800";
    tmp(24942) := x"f800";
    tmp(24943) := x"f800";
    tmp(24944) := x"f800";
    tmp(24945) := x"f800";
    tmp(24946) := x"f800";
    tmp(24947) := x"f800";
    tmp(24948) := x"f800";
    tmp(24949) := x"f800";
    tmp(24950) := x"f800";
    tmp(24951) := x"f800";
    tmp(24952) := x"f800";
    tmp(24953) := x"f800";
    tmp(24954) := x"f800";
    tmp(24955) := x"f800";
    tmp(24956) := x"f800";
    tmp(24957) := x"0840";
    tmp(24958) := x"0840";
    tmp(24959) := x"0840";
    tmp(24960) := x"1040";
    tmp(24961) := x"aa60";
    tmp(24962) := x"9a40";
    tmp(24963) := x"a260";
    tmp(24964) := x"a260";
    tmp(24965) := x"b280";
    tmp(24966) := x"b260";
    tmp(24967) := x"ba80";
    tmp(24968) := x"ca80";
    tmp(24969) := x"cac0";
    tmp(24970) := x"d2c0";
    tmp(24971) := x"dac0";
    tmp(24972) := x"d2a0";
    tmp(24973) := x"d2a0";
    tmp(24974) := x"d2c0";
    tmp(24975) := x"e2e0";
    tmp(24976) := x"e2e0";
    tmp(24977) := x"ca80";
    tmp(24978) := x"c260";
    tmp(24979) := x"c240";
    tmp(24980) := x"ba40";
    tmp(24981) := x"ba60";
    tmp(24982) := x"c280";
    tmp(24983) := x"b260";
    tmp(24984) := x"b260";
    tmp(24985) := x"b240";
    tmp(24986) := x"aa40";
    tmp(24987) := x"aa20";
    tmp(24988) := x"aa20";
    tmp(24989) := x"b240";
    tmp(24990) := x"aa20";
    tmp(24991) := x"b240";
    tmp(24992) := x"aa40";
    tmp(24993) := x"a220";
    tmp(24994) := x"a220";
    tmp(24995) := x"aa60";
    tmp(24996) := x"aa80";
    tmp(24997) := x"b280";
    tmp(24998) := x"aa80";
    tmp(24999) := x"b280";
    tmp(25000) := x"aa60";
    tmp(25001) := x"aa80";
    tmp(25002) := x"aa80";
    tmp(25003) := x"a260";
    tmp(25004) := x"a260";
    tmp(25005) := x"aa60";
    tmp(25006) := x"aa80";
    tmp(25007) := x"b2a0";
    tmp(25008) := x"b2c0";
    tmp(25009) := x"c300";
    tmp(25010) := x"c300";
    tmp(25011) := x"d340";
    tmp(25012) := x"db40";
    tmp(25013) := x"e360";
    tmp(25014) := x"eba0";
    tmp(25015) := x"db60";
    tmp(25016) := x"eba0";
    tmp(25017) := x"ebc0";
    tmp(25018) := x"db80";
    tmp(25019) := x"dba0";
    tmp(25020) := x"cb40";
    tmp(25021) := x"db60";
    tmp(25022) := x"c2c0";
    tmp(25023) := x"baa0";
    tmp(25024) := x"d300";
    tmp(25025) := x"e320";
    tmp(25026) := x"dae0";
    tmp(25027) := x"caa0";
    tmp(25028) := x"d2c0";
    tmp(25029) := x"eb00";
    tmp(25030) := x"fb60";
    tmp(25031) := x"fb80";
    tmp(25032) := x"fb80";
    tmp(25033) := x"eb40";
    tmp(25034) := x"e340";
    tmp(25035) := x"d340";
    tmp(25036) := x"db40";
    tmp(25037) := x"e380";
    tmp(25038) := x"db40";
    tmp(25039) := x"e360";
    tmp(25040) := x"db20";
    tmp(25041) := x"db40";
    tmp(25042) := x"f380";
    tmp(25043) := x"f380";
    tmp(25044) := x"f3a0";
    tmp(25045) := x"f3c0";
    tmp(25046) := x"fba0";
    tmp(25047) := x"fbc0";
    tmp(25048) := x"f360";
    tmp(25049) := x"eb40";
    tmp(25050) := x"eb60";
    tmp(25051) := x"e300";
    tmp(25052) := x"fb80";
    tmp(25053) := x"fb80";
    tmp(25054) := x"e300";
    tmp(25055) := x"79e0";
    tmp(25056) := x"3121";
    tmp(25057) := x"2121";
    tmp(25058) := x"1921";
    tmp(25059) := x"1921";
    tmp(25060) := x"1901";
    tmp(25061) := x"1902";
    tmp(25062) := x"1901";
    tmp(25063) := x"1901";
    tmp(25064) := x"1121";
    tmp(25065) := x"0922";
    tmp(25066) := x"0923";
    tmp(25067) := x"0902";
    tmp(25068) := x"0922";
    tmp(25069) := x"0901";
    tmp(25070) := x"0921";
    tmp(25071) := x"0921";
    tmp(25072) := x"0942";
    tmp(25073) := x"0983";
    tmp(25074) := x"0964";
    tmp(25075) := x"0985";
    tmp(25076) := x"0985";
    tmp(25077) := x"1227";
    tmp(25078) := x"1228";
    tmp(25079) := x"1208";
    tmp(25080) := x"09c8";
    tmp(25081) := x"126a";
    tmp(25082) := x"1b0c";
    tmp(25083) := x"22ca";
    tmp(25084) := x"3b8c";
    tmp(25085) := x"7d10";
    tmp(25086) := x"8c8d";
    tmp(25087) := x"83ea";
    tmp(25088) := x"7baa";
    tmp(25089) := x"6b4a";
    tmp(25090) := x"5b0a";
    tmp(25091) := x"52ea";
    tmp(25092) := x"4288";
    tmp(25093) := x"29e5";
    tmp(25094) := x"2182";
    tmp(25095) := x"1921";
    tmp(25096) := x"2141";
    tmp(25097) := x"29c2";
    tmp(25098) := x"3a23";
    tmp(25099) := x"52a5";
    tmp(25100) := x"6b46";
    tmp(25101) := x"7bc7";
    tmp(25102) := x"9c69";
    tmp(25103) := x"b4eb";
    tmp(25104) := x"c56c";
    tmp(25105) := x"d5ee";
    tmp(25106) := x"e64f";
    tmp(25107) := x"ee8f";
    tmp(25108) := x"ee90";
    tmp(25109) := x"de0f";
    tmp(25110) := x"c56d";
    tmp(25111) := x"bd2d";
    tmp(25112) := x"ac8b";
    tmp(25113) := x"93ea";
    tmp(25114) := x"83a8";
    tmp(25115) := x"7347";
    tmp(25116) := x"6b06";
    tmp(25117) := x"5ac5";
    tmp(25118) := x"5284";
    tmp(25119) := x"4244";
    tmp(25120) := x"4243";
    tmp(25121) := x"4a84";
    tmp(25122) := x"5ac5";
    tmp(25123) := x"6b46";
    tmp(25124) := x"83c8";
    tmp(25125) := x"9c6a";
    tmp(25126) := x"bd2d";
    tmp(25127) := x"d5ef";
    tmp(25128) := x"ee92";
    tmp(25129) := x"ff76";
    tmp(25130) := x"ff98";
    tmp(25131) := x"ffdb";
    tmp(25132) := x"fffe";
    tmp(25133) := x"fffe";
    tmp(25134) := x"fffb";
    tmp(25135) := x"ff98";
    tmp(25136) := x"fef6";
    tmp(25137) := x"e5f3";
    tmp(25138) := x"b4d0";
    tmp(25139) := x"a470";
    tmp(25140) := x"ac91";
    tmp(25141) := x"ac92";
    tmp(25142) := x"b4f3";
    tmp(25143) := x"b4f4";
    tmp(25144) := x"bd15";
    tmp(25145) := x"bd35";
    tmp(25146) := x"c536";
    tmp(25147) := x"b4f5";
    tmp(25148) := x"b515";
    tmp(25149) := x"bcf6";
    tmp(25150) := x"bcf7";
    tmp(25151) := x"bcf7";
    tmp(25152) := x"c537";
    tmp(25153) := x"c537";
    tmp(25154) := x"b4d5";
    tmp(25155) := x"ac95";
    tmp(25156) := x"a475";
    tmp(25157) := x"f800";
    tmp(25158) := x"f800";
    tmp(25159) := x"f800";
    tmp(25160) := x"f800";
    tmp(25161) := x"f800";
    tmp(25162) := x"f800";
    tmp(25163) := x"f800";
    tmp(25164) := x"f800";
    tmp(25165) := x"f800";
    tmp(25166) := x"f800";
    tmp(25167) := x"f800";
    tmp(25168) := x"f800";
    tmp(25169) := x"f800";
    tmp(25170) := x"f800";
    tmp(25171) := x"f800";
    tmp(25172) := x"f800";
    tmp(25173) := x"f800";
    tmp(25174) := x"f800";
    tmp(25175) := x"f800";
    tmp(25176) := x"f800";
    tmp(25177) := x"f800";
    tmp(25178) := x"f800";
    tmp(25179) := x"f800";
    tmp(25180) := x"f800";
    tmp(25181) := x"f800";
    tmp(25182) := x"f800";
    tmp(25183) := x"f800";
    tmp(25184) := x"f800";
    tmp(25185) := x"f800";
    tmp(25186) := x"f800";
    tmp(25187) := x"f800";
    tmp(25188) := x"f800";
    tmp(25189) := x"f800";
    tmp(25190) := x"f800";
    tmp(25191) := x"f800";
    tmp(25192) := x"f800";
    tmp(25193) := x"f800";
    tmp(25194) := x"f800";
    tmp(25195) := x"f800";
    tmp(25196) := x"f800";
    tmp(25197) := x"0840";
    tmp(25198) := x"0840";
    tmp(25199) := x"0840";
    tmp(25200) := x"1040";
    tmp(25201) := x"9a40";
    tmp(25202) := x"9220";
    tmp(25203) := x"9240";
    tmp(25204) := x"9240";
    tmp(25205) := x"a260";
    tmp(25206) := x"aa80";
    tmp(25207) := x"b280";
    tmp(25208) := x"b280";
    tmp(25209) := x"baa0";
    tmp(25210) := x"c2a0";
    tmp(25211) := x"ba80";
    tmp(25212) := x"ba60";
    tmp(25213) := x"b260";
    tmp(25214) := x"c2a0";
    tmp(25215) := x"c2a0";
    tmp(25216) := x"c280";
    tmp(25217) := x"ba60";
    tmp(25218) := x"b220";
    tmp(25219) := x"aa00";
    tmp(25220) := x"aa20";
    tmp(25221) := x"aa20";
    tmp(25222) := x"aa40";
    tmp(25223) := x"aa40";
    tmp(25224) := x"aa40";
    tmp(25225) := x"9a00";
    tmp(25226) := x"9a00";
    tmp(25227) := x"9a00";
    tmp(25228) := x"91c0";
    tmp(25229) := x"91c0";
    tmp(25230) := x"9a00";
    tmp(25231) := x"91c0";
    tmp(25232) := x"89e0";
    tmp(25233) := x"91e0";
    tmp(25234) := x"9200";
    tmp(25235) := x"9220";
    tmp(25236) := x"9220";
    tmp(25237) := x"9200";
    tmp(25238) := x"8a00";
    tmp(25239) := x"8a00";
    tmp(25240) := x"89e0";
    tmp(25241) := x"81c0";
    tmp(25242) := x"81e0";
    tmp(25243) := x"8a00";
    tmp(25244) := x"9a40";
    tmp(25245) := x"9a60";
    tmp(25246) := x"aa80";
    tmp(25247) := x"a280";
    tmp(25248) := x"aaa0";
    tmp(25249) := x"b2e0";
    tmp(25250) := x"cb20";
    tmp(25251) := x"cb20";
    tmp(25252) := x"cb40";
    tmp(25253) := x"db80";
    tmp(25254) := x"db60";
    tmp(25255) := x"d340";
    tmp(25256) := x"c340";
    tmp(25257) := x"c340";
    tmp(25258) := x"c320";
    tmp(25259) := x"dba0";
    tmp(25260) := x"e3c0";
    tmp(25261) := x"9ac0";
    tmp(25262) := x"8200";
    tmp(25263) := x"a280";
    tmp(25264) := x"c2e0";
    tmp(25265) := x"d300";
    tmp(25266) := x"d2e0";
    tmp(25267) := x"d2c0";
    tmp(25268) := x"dac0";
    tmp(25269) := x"eb20";
    tmp(25270) := x"f340";
    tmp(25271) := x"fb80";
    tmp(25272) := x"e340";
    tmp(25273) := x"bae0";
    tmp(25274) := x"aaa0";
    tmp(25275) := x"9a80";
    tmp(25276) := x"a2c0";
    tmp(25277) := x"aac0";
    tmp(25278) := x"aac0";
    tmp(25279) := x"b2c0";
    tmp(25280) := x"bae0";
    tmp(25281) := x"c320";
    tmp(25282) := x"cb40";
    tmp(25283) := x"cb20";
    tmp(25284) := x"db40";
    tmp(25285) := x"db40";
    tmp(25286) := x"eb60";
    tmp(25287) := x"e360";
    tmp(25288) := x"e360";
    tmp(25289) := x"db20";
    tmp(25290) := x"d300";
    tmp(25291) := x"db40";
    tmp(25292) := x"f380";
    tmp(25293) := x"f360";
    tmp(25294) := x"b2a0";
    tmp(25295) := x"4980";
    tmp(25296) := x"2122";
    tmp(25297) := x"1123";
    tmp(25298) := x"1123";
    tmp(25299) := x"1123";
    tmp(25300) := x"1124";
    tmp(25301) := x"1104";
    tmp(25302) := x"1123";
    tmp(25303) := x"0902";
    tmp(25304) := x"08e2";
    tmp(25305) := x"0902";
    tmp(25306) := x"0902";
    tmp(25307) := x"0901";
    tmp(25308) := x"0942";
    tmp(25309) := x"0942";
    tmp(25310) := x"0922";
    tmp(25311) := x"0942";
    tmp(25312) := x"0983";
    tmp(25313) := x"11a4";
    tmp(25314) := x"11c5";
    tmp(25315) := x"1207";
    tmp(25316) := x"1207";
    tmp(25317) := x"11c7";
    tmp(25318) := x"11e8";
    tmp(25319) := x"09e8";
    tmp(25320) := x"128a";
    tmp(25321) := x"232a";
    tmp(25322) := x"3369";
    tmp(25323) := x"4b68";
    tmp(25324) := x"740a";
    tmp(25325) := x"8c0a";
    tmp(25326) := x"944b";
    tmp(25327) := x"944b";
    tmp(25328) := x"83eb";
    tmp(25329) := x"73ac";
    tmp(25330) := x"6b6c";
    tmp(25331) := x"634c";
    tmp(25332) := x"52eb";
    tmp(25333) := x"3a67";
    tmp(25334) := x"29a3";
    tmp(25335) := x"1942";
    tmp(25336) := x"1921";
    tmp(25337) := x"1941";
    tmp(25338) := x"29a2";
    tmp(25339) := x"3a03";
    tmp(25340) := x"4a84";
    tmp(25341) := x"6325";
    tmp(25342) := x"7bc7";
    tmp(25343) := x"9448";
    tmp(25344) := x"acca";
    tmp(25345) := x"c58d";
    tmp(25346) := x"de0f";
    tmp(25347) := x"e62f";
    tmp(25348) := x"ee90";
    tmp(25349) := x"e64f";
    tmp(25350) := x"e60f";
    tmp(25351) := x"cd6e";
    tmp(25352) := x"bced";
    tmp(25353) := x"ac8b";
    tmp(25354) := x"940a";
    tmp(25355) := x"8bc9";
    tmp(25356) := x"7367";
    tmp(25357) := x"6b26";
    tmp(25358) := x"5ac5";
    tmp(25359) := x"52a5";
    tmp(25360) := x"4244";
    tmp(25361) := x"4243";
    tmp(25362) := x"4a64";
    tmp(25363) := x"5ac5";
    tmp(25364) := x"6b46";
    tmp(25365) := x"7ba8";
    tmp(25366) := x"9c6a";
    tmp(25367) := x"ad0d";
    tmp(25368) := x"cdaf";
    tmp(25369) := x"ee73";
    tmp(25370) := x"fef5";
    tmp(25371) := x"ff78";
    tmp(25372) := x"ffda";
    tmp(25373) := x"ffba";
    tmp(25374) := x"ffdb";
    tmp(25375) := x"ff78";
    tmp(25376) := x"ff16";
    tmp(25377) := x"ddd3";
    tmp(25378) := x"bcf1";
    tmp(25379) := x"ac91";
    tmp(25380) := x"acb1";
    tmp(25381) := x"bcf3";
    tmp(25382) := x"bcf4";
    tmp(25383) := x"bd15";
    tmp(25384) := x"bd35";
    tmp(25385) := x"bd35";
    tmp(25386) := x"bd76";
    tmp(25387) := x"bd35";
    tmp(25388) := x"bd15";
    tmp(25389) := x"bd16";
    tmp(25390) := x"bd17";
    tmp(25391) := x"c517";
    tmp(25392) := x"bcf6";
    tmp(25393) := x"bd36";
    tmp(25394) := x"bcf6";
    tmp(25395) := x"ac95";
    tmp(25396) := x"ac95";
    tmp(25397) := x"f800";
    tmp(25398) := x"f800";
    tmp(25399) := x"f800";
    tmp(25400) := x"f800";
    tmp(25401) := x"f800";
    tmp(25402) := x"f800";
    tmp(25403) := x"f800";
    tmp(25404) := x"f800";
    tmp(25405) := x"f800";
    tmp(25406) := x"f800";
    tmp(25407) := x"f800";
    tmp(25408) := x"f800";
    tmp(25409) := x"f800";
    tmp(25410) := x"f800";
    tmp(25411) := x"f800";
    tmp(25412) := x"f800";
    tmp(25413) := x"f800";
    tmp(25414) := x"f800";
    tmp(25415) := x"f800";
    tmp(25416) := x"f800";
    tmp(25417) := x"f800";
    tmp(25418) := x"f800";
    tmp(25419) := x"f800";
    tmp(25420) := x"f800";
    tmp(25421) := x"f800";
    tmp(25422) := x"f800";
    tmp(25423) := x"f800";
    tmp(25424) := x"f800";
    tmp(25425) := x"f800";
    tmp(25426) := x"f800";
    tmp(25427) := x"f800";
    tmp(25428) := x"f800";
    tmp(25429) := x"f800";
    tmp(25430) := x"f800";
    tmp(25431) := x"f800";
    tmp(25432) := x"f800";
    tmp(25433) := x"f800";
    tmp(25434) := x"f800";
    tmp(25435) := x"f800";
    tmp(25436) := x"f800";
    tmp(25437) := x"0840";
    tmp(25438) := x"0840";
    tmp(25439) := x"0840";
    tmp(25440) := x"1040";
    tmp(25441) := x"9240";
    tmp(25442) := x"8220";
    tmp(25443) := x"8a40";
    tmp(25444) := x"8a40";
    tmp(25445) := x"9aa0";
    tmp(25446) := x"b300";
    tmp(25447) := x"b300";
    tmp(25448) := x"b2e0";
    tmp(25449) := x"aaa0";
    tmp(25450) := x"b280";
    tmp(25451) := x"aa60";
    tmp(25452) := x"9a20";
    tmp(25453) := x"9220";
    tmp(25454) := x"9a20";
    tmp(25455) := x"a260";
    tmp(25456) := x"a240";
    tmp(25457) := x"a220";
    tmp(25458) := x"9a00";
    tmp(25459) := x"91e0";
    tmp(25460) := x"91e0";
    tmp(25461) := x"91e0";
    tmp(25462) := x"99e0";
    tmp(25463) := x"91e0";
    tmp(25464) := x"91e0";
    tmp(25465) := x"89e0";
    tmp(25466) := x"89c0";
    tmp(25467) := x"81a0";
    tmp(25468) := x"81a0";
    tmp(25469) := x"81a0";
    tmp(25470) := x"81a0";
    tmp(25471) := x"7980";
    tmp(25472) := x"79a0";
    tmp(25473) := x"79a0";
    tmp(25474) := x"79a0";
    tmp(25475) := x"79a0";
    tmp(25476) := x"79c0";
    tmp(25477) := x"79a0";
    tmp(25478) := x"71a0";
    tmp(25479) := x"71a0";
    tmp(25480) := x"6960";
    tmp(25481) := x"6140";
    tmp(25482) := x"6160";
    tmp(25483) := x"6980";
    tmp(25484) := x"79c0";
    tmp(25485) := x"8a00";
    tmp(25486) := x"9a40";
    tmp(25487) := x"9a40";
    tmp(25488) := x"b2c0";
    tmp(25489) := x"aac0";
    tmp(25490) := x"bae0";
    tmp(25491) := x"bb00";
    tmp(25492) := x"c340";
    tmp(25493) := x"bb20";
    tmp(25494) := x"bb00";
    tmp(25495) := x"aae0";
    tmp(25496) := x"aac0";
    tmp(25497) := x"b300";
    tmp(25498) := x"bb20";
    tmp(25499) := x"b340";
    tmp(25500) := x"82a0";
    tmp(25501) := x"3920";
    tmp(25502) := x"59a0";
    tmp(25503) := x"8a60";
    tmp(25504) := x"a2a0";
    tmp(25505) := x"aa80";
    tmp(25506) := x"c2c0";
    tmp(25507) := x"db20";
    tmp(25508) := x"e320";
    tmp(25509) := x"eb20";
    tmp(25510) := x"f360";
    tmp(25511) := x"fb80";
    tmp(25512) := x"c2e0";
    tmp(25513) := x"8240";
    tmp(25514) := x"6a20";
    tmp(25515) := x"51e0";
    tmp(25516) := x"5a00";
    tmp(25517) := x"6a20";
    tmp(25518) := x"7a40";
    tmp(25519) := x"8a60";
    tmp(25520) := x"92a0";
    tmp(25521) := x"9aa0";
    tmp(25522) := x"9a80";
    tmp(25523) := x"9a80";
    tmp(25524) := x"aac0";
    tmp(25525) := x"b2c0";
    tmp(25526) := x"b2c0";
    tmp(25527) := x"b2c0";
    tmp(25528) := x"aac0";
    tmp(25529) := x"b2c0";
    tmp(25530) := x"cb20";
    tmp(25531) := x"d320";
    tmp(25532) := x"db20";
    tmp(25533) := x"c320";
    tmp(25534) := x"6200";
    tmp(25535) := x"2161";
    tmp(25536) := x"1163";
    tmp(25537) := x"1144";
    tmp(25538) := x"0924";
    tmp(25539) := x"0924";
    tmp(25540) := x"1145";
    tmp(25541) := x"1165";
    tmp(25542) := x"0925";
    tmp(25543) := x"08e3";
    tmp(25544) := x"0903";
    tmp(25545) := x"0943";
    tmp(25546) := x"0902";
    tmp(25547) := x"0922";
    tmp(25548) := x"0984";
    tmp(25549) := x"0985";
    tmp(25550) := x"11c6";
    tmp(25551) := x"11e6";
    tmp(25552) := x"11c6";
    tmp(25553) := x"11c5";
    tmp(25554) := x"11e7";
    tmp(25555) := x"1248";
    tmp(25556) := x"1208";
    tmp(25557) := x"0945";
    tmp(25558) := x"1185";
    tmp(25559) := x"19e5";
    tmp(25560) := x"1a04";
    tmp(25561) := x"19c2";
    tmp(25562) := x"2a02";
    tmp(25563) := x"4283";
    tmp(25564) := x"5b06";
    tmp(25565) := x"7bc8";
    tmp(25566) := x"8c4a";
    tmp(25567) := x"944b";
    tmp(25568) := x"8c0c";
    tmp(25569) := x"83ed";
    tmp(25570) := x"7bee";
    tmp(25571) := x"73ce";
    tmp(25572) := x"634d";
    tmp(25573) := x"4ac9";
    tmp(25574) := x"3205";
    tmp(25575) := x"2182";
    tmp(25576) := x"1941";
    tmp(25577) := x"1921";
    tmp(25578) := x"1941";
    tmp(25579) := x"29a2";
    tmp(25580) := x"3202";
    tmp(25581) := x"4a84";
    tmp(25582) := x"6325";
    tmp(25583) := x"7b86";
    tmp(25584) := x"9408";
    tmp(25585) := x"acaa";
    tmp(25586) := x"bd4c";
    tmp(25587) := x"cdae";
    tmp(25588) := x"e670";
    tmp(25589) := x"ee90";
    tmp(25590) := x"ee50";
    tmp(25591) := x"ddef";
    tmp(25592) := x"c56e";
    tmp(25593) := x"b4ec";
    tmp(25594) := x"a48b";
    tmp(25595) := x"9c2a";
    tmp(25596) := x"83a9";
    tmp(25597) := x"7367";
    tmp(25598) := x"6b26";
    tmp(25599) := x"5ae6";
    tmp(25600) := x"52a5";
    tmp(25601) := x"4a64";
    tmp(25602) := x"4244";
    tmp(25603) := x"4a64";
    tmp(25604) := x"5ac5";
    tmp(25605) := x"6b26";
    tmp(25606) := x"7ba8";
    tmp(25607) := x"946a";
    tmp(25608) := x"accc";
    tmp(25609) := x"c58f";
    tmp(25610) := x"e612";
    tmp(25611) := x"ee94";
    tmp(25612) := x"ff16";
    tmp(25613) := x"ff57";
    tmp(25614) := x"ff78";
    tmp(25615) := x"ff58";
    tmp(25616) := x"f6b6";
    tmp(25617) := x"d5d2";
    tmp(25618) := x"b4f1";
    tmp(25619) := x"b4f2";
    tmp(25620) := x"b4f3";
    tmp(25621) := x"bd34";
    tmp(25622) := x"bd34";
    tmp(25623) := x"c575";
    tmp(25624) := x"bd35";
    tmp(25625) := x"bd56";
    tmp(25626) := x"c576";
    tmp(25627) := x"bd56";
    tmp(25628) := x"bd36";
    tmp(25629) := x"bd36";
    tmp(25630) := x"bd37";
    tmp(25631) := x"bd17";
    tmp(25632) := x"c556";
    tmp(25633) := x"bcf6";
    tmp(25634) := x"b4d5";
    tmp(25635) := x"a494";
    tmp(25636) := x"ac94";
    tmp(25637) := x"f800";
    tmp(25638) := x"f800";
    tmp(25639) := x"f800";
    tmp(25640) := x"f800";
    tmp(25641) := x"f800";
    tmp(25642) := x"f800";
    tmp(25643) := x"f800";
    tmp(25644) := x"f800";
    tmp(25645) := x"f800";
    tmp(25646) := x"f800";
    tmp(25647) := x"f800";
    tmp(25648) := x"f800";
    tmp(25649) := x"f800";
    tmp(25650) := x"f800";
    tmp(25651) := x"f800";
    tmp(25652) := x"f800";
    tmp(25653) := x"f800";
    tmp(25654) := x"f800";
    tmp(25655) := x"f800";
    tmp(25656) := x"f800";
    tmp(25657) := x"f800";
    tmp(25658) := x"f800";
    tmp(25659) := x"f800";
    tmp(25660) := x"f800";
    tmp(25661) := x"f800";
    tmp(25662) := x"f800";
    tmp(25663) := x"f800";
    tmp(25664) := x"f800";
    tmp(25665) := x"f800";
    tmp(25666) := x"f800";
    tmp(25667) := x"f800";
    tmp(25668) := x"f800";
    tmp(25669) := x"f800";
    tmp(25670) := x"f800";
    tmp(25671) := x"f800";
    tmp(25672) := x"f800";
    tmp(25673) := x"f800";
    tmp(25674) := x"f800";
    tmp(25675) := x"f800";
    tmp(25676) := x"f800";
    tmp(25677) := x"0840";
    tmp(25678) := x"0840";
    tmp(25679) := x"0840";
    tmp(25680) := x"0820";
    tmp(25681) := x"79e0";
    tmp(25682) := x"7200";
    tmp(25683) := x"7a00";
    tmp(25684) := x"7a20";
    tmp(25685) := x"7a40";
    tmp(25686) := x"7a40";
    tmp(25687) := x"8240";
    tmp(25688) := x"8a60";
    tmp(25689) := x"9240";
    tmp(25690) := x"9220";
    tmp(25691) := x"8a00";
    tmp(25692) := x"8a00";
    tmp(25693) := x"81e0";
    tmp(25694) := x"8a00";
    tmp(25695) := x"89e0";
    tmp(25696) := x"91e0";
    tmp(25697) := x"89c0";
    tmp(25698) := x"89a0";
    tmp(25699) := x"81a0";
    tmp(25700) := x"81a0";
    tmp(25701) := x"8180";
    tmp(25702) := x"81a0";
    tmp(25703) := x"7980";
    tmp(25704) := x"7980";
    tmp(25705) := x"7980";
    tmp(25706) := x"7980";
    tmp(25707) := x"7180";
    tmp(25708) := x"7160";
    tmp(25709) := x"7160";
    tmp(25710) := x"6960";
    tmp(25711) := x"6940";
    tmp(25712) := x"6140";
    tmp(25713) := x"6940";
    tmp(25714) := x"6140";
    tmp(25715) := x"5940";
    tmp(25716) := x"5940";
    tmp(25717) := x"5940";
    tmp(25718) := x"5140";
    tmp(25719) := x"5140";
    tmp(25720) := x"4120";
    tmp(25721) := x"3900";
    tmp(25722) := x"3900";
    tmp(25723) := x"3900";
    tmp(25724) := x"4980";
    tmp(25725) := x"59c0";
    tmp(25726) := x"71e0";
    tmp(25727) := x"8220";
    tmp(25728) := x"8a40";
    tmp(25729) := x"9aa0";
    tmp(25730) := x"aac0";
    tmp(25731) := x"b300";
    tmp(25732) := x"bb20";
    tmp(25733) := x"aac0";
    tmp(25734) := x"a2a0";
    tmp(25735) := x"9a80";
    tmp(25736) := x"9280";
    tmp(25737) := x"9280";
    tmp(25738) := x"9ae0";
    tmp(25739) := x"6a60";
    tmp(25740) := x"18e1";
    tmp(25741) := x"20e0";
    tmp(25742) := x"4180";
    tmp(25743) := x"51a0";
    tmp(25744) := x"69e0";
    tmp(25745) := x"8a60";
    tmp(25746) := x"aac0";
    tmp(25747) := x"c2e0";
    tmp(25748) := x"c2c0";
    tmp(25749) := x"db00";
    tmp(25750) := x"f360";
    tmp(25751) := x"f360";
    tmp(25752) := x"b2c0";
    tmp(25753) := x"7241";
    tmp(25754) := x"41e2";
    tmp(25755) := x"2962";
    tmp(25756) := x"39a1";
    tmp(25757) := x"41a0";
    tmp(25758) := x"49a0";
    tmp(25759) := x"59e0";
    tmp(25760) := x"6a40";
    tmp(25761) := x"6a20";
    tmp(25762) := x"6200";
    tmp(25763) := x"6a20";
    tmp(25764) := x"7220";
    tmp(25765) := x"7240";
    tmp(25766) := x"6a20";
    tmp(25767) := x"6a00";
    tmp(25768) := x"6a00";
    tmp(25769) := x"8a60";
    tmp(25770) := x"a2c0";
    tmp(25771) := x"a280";
    tmp(25772) := x"aac0";
    tmp(25773) := x"7280";
    tmp(25774) := x"29a1";
    tmp(25775) := x"1184";
    tmp(25776) := x"11a5";
    tmp(25777) := x"0965";
    tmp(25778) := x"0945";
    tmp(25779) := x"0945";
    tmp(25780) := x"1186";
    tmp(25781) := x"1186";
    tmp(25782) := x"0924";
    tmp(25783) := x"0904";
    tmp(25784) := x"0924";
    tmp(25785) := x"0965";
    tmp(25786) := x"0985";
    tmp(25787) := x"11a5";
    tmp(25788) := x"1185";
    tmp(25789) := x"11a6";
    tmp(25790) := x"11c6";
    tmp(25791) := x"11c6";
    tmp(25792) := x"1a07";
    tmp(25793) := x"2aca";
    tmp(25794) := x"32ea";
    tmp(25795) := x"32a9";
    tmp(25796) := x"32c9";
    tmp(25797) := x"3a87";
    tmp(25798) := x"3a85";
    tmp(25799) := x"2a02";
    tmp(25800) := x"1961";
    tmp(25801) := x"1120";
    tmp(25802) := x"1981";
    tmp(25803) := x"3202";
    tmp(25804) := x"4aa4";
    tmp(25805) := x"6346";
    tmp(25806) := x"7be9";
    tmp(25807) := x"944a";
    tmp(25808) := x"944b";
    tmp(25809) := x"944d";
    tmp(25810) := x"8c6f";
    tmp(25811) := x"7c10";
    tmp(25812) := x"6bcf";
    tmp(25813) := x"5b4b";
    tmp(25814) := x"4287";
    tmp(25815) := x"31e3";
    tmp(25816) := x"2162";
    tmp(25817) := x"1921";
    tmp(25818) := x"1921";
    tmp(25819) := x"1941";
    tmp(25820) := x"2181";
    tmp(25821) := x"3202";
    tmp(25822) := x"4a83";
    tmp(25823) := x"5ae5";
    tmp(25824) := x"7366";
    tmp(25825) := x"8be8";
    tmp(25826) := x"a4aa";
    tmp(25827) := x"b52b";
    tmp(25828) := x"d5ed";
    tmp(25829) := x"ee2f";
    tmp(25830) := x"ee91";
    tmp(25831) := x"ee50";
    tmp(25832) := x"d5cf";
    tmp(25833) := x"cd6e";
    tmp(25834) := x"bced";
    tmp(25835) := x"ac8b";
    tmp(25836) := x"940a";
    tmp(25837) := x"83a8";
    tmp(25838) := x"7367";
    tmp(25839) := x"6b27";
    tmp(25840) := x"62e6";
    tmp(25841) := x"52a5";
    tmp(25842) := x"4a64";
    tmp(25843) := x"4a64";
    tmp(25844) := x"4a64";
    tmp(25845) := x"52a5";
    tmp(25846) := x"6326";
    tmp(25847) := x"7b88";
    tmp(25848) := x"940a";
    tmp(25849) := x"a48c";
    tmp(25850) := x"bd2f";
    tmp(25851) := x"cdb0";
    tmp(25852) := x"e632";
    tmp(25853) := x"ee95";
    tmp(25854) := x"f6d6";
    tmp(25855) := x"feb6";
    tmp(25856) := x"ee95";
    tmp(25857) := x"cdb3";
    tmp(25858) := x"bd12";
    tmp(25859) := x"b4f2";
    tmp(25860) := x"bd13";
    tmp(25861) := x"bd34";
    tmp(25862) := x"c575";
    tmp(25863) := x"c5b6";
    tmp(25864) := x"c576";
    tmp(25865) := x"bd56";
    tmp(25866) := x"c5b7";
    tmp(25867) := x"c576";
    tmp(25868) := x"c535";
    tmp(25869) := x"bd16";
    tmp(25870) := x"c558";
    tmp(25871) := x"bd17";
    tmp(25872) := x"c536";
    tmp(25873) := x"bd16";
    tmp(25874) := x"bcd6";
    tmp(25875) := x"b4b5";
    tmp(25876) := x"b4b5";
    tmp(25877) := x"f800";
    tmp(25878) := x"f800";
    tmp(25879) := x"f800";
    tmp(25880) := x"f800";
    tmp(25881) := x"f800";
    tmp(25882) := x"f800";
    tmp(25883) := x"f800";
    tmp(25884) := x"f800";
    tmp(25885) := x"f800";
    tmp(25886) := x"f800";
    tmp(25887) := x"f800";
    tmp(25888) := x"f800";
    tmp(25889) := x"f800";
    tmp(25890) := x"f800";
    tmp(25891) := x"f800";
    tmp(25892) := x"f800";
    tmp(25893) := x"f800";
    tmp(25894) := x"f800";
    tmp(25895) := x"f800";
    tmp(25896) := x"f800";
    tmp(25897) := x"f800";
    tmp(25898) := x"f800";
    tmp(25899) := x"f800";
    tmp(25900) := x"f800";
    tmp(25901) := x"f800";
    tmp(25902) := x"f800";
    tmp(25903) := x"f800";
    tmp(25904) := x"f800";
    tmp(25905) := x"f800";
    tmp(25906) := x"f800";
    tmp(25907) := x"f800";
    tmp(25908) := x"f800";
    tmp(25909) := x"f800";
    tmp(25910) := x"f800";
    tmp(25911) := x"f800";
    tmp(25912) := x"f800";
    tmp(25913) := x"f800";
    tmp(25914) := x"f800";
    tmp(25915) := x"f800";
    tmp(25916) := x"f800";
    tmp(25917) := x"0840";
    tmp(25918) := x"0840";
    tmp(25919) := x"0840";
    tmp(25920) := x"0820";
    tmp(25921) := x"69c0";
    tmp(25922) := x"61a0";
    tmp(25923) := x"61a0";
    tmp(25924) := x"61c0";
    tmp(25925) := x"59c0";
    tmp(25926) := x"59c0";
    tmp(25927) := x"61a0";
    tmp(25928) := x"6180";
    tmp(25929) := x"6180";
    tmp(25930) := x"6180";
    tmp(25931) := x"6180";
    tmp(25932) := x"5960";
    tmp(25933) := x"6180";
    tmp(25934) := x"6980";
    tmp(25935) := x"6160";
    tmp(25936) := x"6980";
    tmp(25937) := x"6960";
    tmp(25938) := x"6940";
    tmp(25939) := x"6940";
    tmp(25940) := x"6940";
    tmp(25941) := x"6940";
    tmp(25942) := x"6940";
    tmp(25943) := x"6120";
    tmp(25944) := x"6120";
    tmp(25945) := x"5900";
    tmp(25946) := x"5920";
    tmp(25947) := x"5920";
    tmp(25948) := x"5100";
    tmp(25949) := x"5100";
    tmp(25950) := x"4900";
    tmp(25951) := x"4900";
    tmp(25952) := x"4920";
    tmp(25953) := x"4940";
    tmp(25954) := x"4140";
    tmp(25955) := x"4140";
    tmp(25956) := x"3120";
    tmp(25957) := x"3140";
    tmp(25958) := x"2961";
    tmp(25959) := x"2141";
    tmp(25960) := x"1901";
    tmp(25961) := x"10e1";
    tmp(25962) := x"10c1";
    tmp(25963) := x"10c1";
    tmp(25964) := x"1963";
    tmp(25965) := x"1982";
    tmp(25966) := x"2161";
    tmp(25967) := x"39c1";
    tmp(25968) := x"5200";
    tmp(25969) := x"6a20";
    tmp(25970) := x"7a40";
    tmp(25971) := x"9aa0";
    tmp(25972) := x"9ac0";
    tmp(25973) := x"9aa0";
    tmp(25974) := x"8a60";
    tmp(25975) := x"7a20";
    tmp(25976) := x"6a20";
    tmp(25977) := x"6a40";
    tmp(25978) := x"5221";
    tmp(25979) := x"1941";
    tmp(25980) := x"08a1";
    tmp(25981) := x"10e1";
    tmp(25982) := x"18e0";
    tmp(25983) := x"2900";
    tmp(25984) := x"51a0";
    tmp(25985) := x"7a40";
    tmp(25986) := x"9280";
    tmp(25987) := x"9a80";
    tmp(25988) := x"aaa0";
    tmp(25989) := x"cb00";
    tmp(25990) := x"db20";
    tmp(25991) := x"eb60";
    tmp(25992) := x"cb20";
    tmp(25993) := x"8281";
    tmp(25994) := x"2983";
    tmp(25995) := x"1943";
    tmp(25996) := x"1942";
    tmp(25997) := x"2982";
    tmp(25998) := x"29a1";
    tmp(25999) := x"31a1";
    tmp(26000) := x"3181";
    tmp(26001) := x"3181";
    tmp(26002) := x"3160";
    tmp(26003) := x"3180";
    tmp(26004) := x"3181";
    tmp(26005) := x"39a1";
    tmp(26006) := x"39a1";
    tmp(26007) := x"3980";
    tmp(26008) := x"49a0";
    tmp(26009) := x"5a00";
    tmp(26010) := x"6240";
    tmp(26011) := x"6240";
    tmp(26012) := x"4a01";
    tmp(26013) := x"2161";
    tmp(26014) := x"1143";
    tmp(26015) := x"1165";
    tmp(26016) := x"11a6";
    tmp(26017) := x"0945";
    tmp(26018) := x"0945";
    tmp(26019) := x"1186";
    tmp(26020) := x"11a6";
    tmp(26021) := x"0945";
    tmp(26022) := x"0904";
    tmp(26023) := x"0924";
    tmp(26024) := x"0965";
    tmp(26025) := x"11c6";
    tmp(26026) := x"11e7";
    tmp(26027) := x"11a7";
    tmp(26028) := x"1166";
    tmp(26029) := x"19e7";
    tmp(26030) := x"3b2c";
    tmp(26031) := x"5c0f";
    tmp(26032) := x"7cf2";
    tmp(26033) := x"9e15";
    tmp(26034) := x"9db2";
    tmp(26035) := x"956f";
    tmp(26036) := x"9daf";
    tmp(26037) := x"7c8a";
    tmp(26038) := x"5345";
    tmp(26039) := x"2a22";
    tmp(26040) := x"1140";
    tmp(26041) := x"08e0";
    tmp(26042) := x"1120";
    tmp(26043) := x"21a1";
    tmp(26044) := x"3a43";
    tmp(26045) := x"52c5";
    tmp(26046) := x"6b67";
    tmp(26047) := x"83e8";
    tmp(26048) := x"8c4a";
    tmp(26049) := x"946d";
    tmp(26050) := x"94b1";
    tmp(26051) := x"8c72";
    tmp(26052) := x"8451";
    tmp(26053) := x"6b8d";
    tmp(26054) := x"52e9";
    tmp(26055) := x"3a25";
    tmp(26056) := x"29a3";
    tmp(26057) := x"1941";
    tmp(26058) := x"1921";
    tmp(26059) := x"1121";
    tmp(26060) := x"1921";
    tmp(26061) := x"2181";
    tmp(26062) := x"31e2";
    tmp(26063) := x"4263";
    tmp(26064) := x"5ac4";
    tmp(26065) := x"7346";
    tmp(26066) := x"8be7";
    tmp(26067) := x"9c89";
    tmp(26068) := x"bd4b";
    tmp(26069) := x"cd8d";
    tmp(26070) := x"ddef";
    tmp(26071) := x"ee50";
    tmp(26072) := x"e630";
    tmp(26073) := x"e610";
    tmp(26074) := x"cd6e";
    tmp(26075) := x"bced";
    tmp(26076) := x"ac6b";
    tmp(26077) := x"93ea";
    tmp(26078) := x"83a8";
    tmp(26079) := x"7368";
    tmp(26080) := x"6b27";
    tmp(26081) := x"62e6";
    tmp(26082) := x"52a5";
    tmp(26083) := x"4a84";
    tmp(26084) := x"4a64";
    tmp(26085) := x"4a85";
    tmp(26086) := x"5285";
    tmp(26087) := x"6b06";
    tmp(26088) := x"7b68";
    tmp(26089) := x"8bea";
    tmp(26090) := x"a46c";
    tmp(26091) := x"b4ee";
    tmp(26092) := x"c550";
    tmp(26093) := x"cdd2";
    tmp(26094) := x"ddf4";
    tmp(26095) := x"e634";
    tmp(26096) := x"de34";
    tmp(26097) := x"c572";
    tmp(26098) := x"c553";
    tmp(26099) := x"bd13";
    tmp(26100) := x"bcf3";
    tmp(26101) := x"bd14";
    tmp(26102) := x"c595";
    tmp(26103) := x"cdb6";
    tmp(26104) := x"c597";
    tmp(26105) := x"c576";
    tmp(26106) := x"c577";
    tmp(26107) := x"c597";
    tmp(26108) := x"c577";
    tmp(26109) := x"c537";
    tmp(26110) := x"c537";
    tmp(26111) := x"bd17";
    tmp(26112) := x"c536";
    tmp(26113) := x"bcf5";
    tmp(26114) := x"b4d6";
    tmp(26115) := x"ac95";
    tmp(26116) := x"b4b6";
    tmp(26117) := x"f800";
    tmp(26118) := x"f800";
    tmp(26119) := x"f800";
    tmp(26120) := x"f800";
    tmp(26121) := x"f800";
    tmp(26122) := x"f800";
    tmp(26123) := x"f800";
    tmp(26124) := x"f800";
    tmp(26125) := x"f800";
    tmp(26126) := x"f800";
    tmp(26127) := x"f800";
    tmp(26128) := x"f800";
    tmp(26129) := x"f800";
    tmp(26130) := x"f800";
    tmp(26131) := x"f800";
    tmp(26132) := x"f800";
    tmp(26133) := x"f800";
    tmp(26134) := x"f800";
    tmp(26135) := x"f800";
    tmp(26136) := x"f800";
    tmp(26137) := x"f800";
    tmp(26138) := x"f800";
    tmp(26139) := x"f800";
    tmp(26140) := x"f800";
    tmp(26141) := x"f800";
    tmp(26142) := x"f800";
    tmp(26143) := x"f800";
    tmp(26144) := x"f800";
    tmp(26145) := x"f800";
    tmp(26146) := x"f800";
    tmp(26147) := x"f800";
    tmp(26148) := x"f800";
    tmp(26149) := x"f800";
    tmp(26150) := x"f800";
    tmp(26151) := x"f800";
    tmp(26152) := x"f800";
    tmp(26153) := x"f800";
    tmp(26154) := x"f800";
    tmp(26155) := x"f800";
    tmp(26156) := x"f800";
    tmp(26157) := x"0840";
    tmp(26158) := x"0840";
    tmp(26159) := x"0840";
    tmp(26160) := x"0820";
    tmp(26161) := x"4960";
    tmp(26162) := x"4140";
    tmp(26163) := x"4160";
    tmp(26164) := x"4160";
    tmp(26165) := x"3940";
    tmp(26166) := x"3100";
    tmp(26167) := x"30e0";
    tmp(26168) := x"3100";
    tmp(26169) := x"3900";
    tmp(26170) := x"4120";
    tmp(26171) := x"61e1";
    tmp(26172) := x"6a41";
    tmp(26173) := x"6a21";
    tmp(26174) := x"51a0";
    tmp(26175) := x"4160";
    tmp(26176) := x"4120";
    tmp(26177) := x"5980";
    tmp(26178) := x"61c0";
    tmp(26179) := x"51a0";
    tmp(26180) := x"5180";
    tmp(26181) := x"4960";
    tmp(26182) := x"4960";
    tmp(26183) := x"4920";
    tmp(26184) := x"4100";
    tmp(26185) := x"4140";
    tmp(26186) := x"3940";
    tmp(26187) := x"3140";
    tmp(26188) := x"3961";
    tmp(26189) := x"3161";
    tmp(26190) := x"39a1";
    tmp(26191) := x"2961";
    tmp(26192) := x"1921";
    tmp(26193) := x"1962";
    tmp(26194) := x"1122";
    tmp(26195) := x"1102";
    tmp(26196) := x"08c2";
    tmp(26197) := x"0903";
    tmp(26198) := x"0924";
    tmp(26199) := x"0904";
    tmp(26200) := x"0904";
    tmp(26201) := x"0905";
    tmp(26202) := x"1145";
    tmp(26203) := x"0904";
    tmp(26204) := x"0925";
    tmp(26205) := x"0946";
    tmp(26206) := x"0925";
    tmp(26207) := x"1145";
    tmp(26208) := x"1964";
    tmp(26209) := x"2162";
    tmp(26210) := x"39a1";
    tmp(26211) := x"51c0";
    tmp(26212) := x"7240";
    tmp(26213) := x"7a40";
    tmp(26214) := x"6a00";
    tmp(26215) := x"51e1";
    tmp(26216) := x"39a1";
    tmp(26217) := x"2981";
    tmp(26218) := x"1122";
    tmp(26219) := x"08c3";
    tmp(26220) := x"08c3";
    tmp(26221) := x"08a2";
    tmp(26222) := x"08a1";
    tmp(26223) := x"2100";
    tmp(26224) := x"41a0";
    tmp(26225) := x"6200";
    tmp(26226) := x"7240";
    tmp(26227) := x"8a80";
    tmp(26228) := x"9aa0";
    tmp(26229) := x"b2e0";
    tmp(26230) := x"c300";
    tmp(26231) := x"cb40";
    tmp(26232) := x"bae0";
    tmp(26233) := x"7241";
    tmp(26234) := x"2163";
    tmp(26235) := x"1103";
    tmp(26236) := x"1124";
    tmp(26237) := x"1124";
    tmp(26238) := x"1164";
    tmp(26239) := x"1963";
    tmp(26240) := x"1122";
    tmp(26241) := x"1102";
    tmp(26242) := x"1102";
    tmp(26243) := x"1122";
    tmp(26244) := x"1122";
    tmp(26245) := x"1962";
    tmp(26246) := x"2183";
    tmp(26247) := x"2982";
    tmp(26248) := x"29c2";
    tmp(26249) := x"29a2";
    tmp(26250) := x"2182";
    tmp(26251) := x"1982";
    tmp(26252) := x"1123";
    tmp(26253) := x"0944";
    tmp(26254) := x"1185";
    tmp(26255) := x"1186";
    tmp(26256) := x"0965";
    tmp(26257) := x"0965";
    tmp(26258) := x"0986";
    tmp(26259) := x"1187";
    tmp(26260) := x"11a7";
    tmp(26261) := x"11a7";
    tmp(26262) := x"09a7";
    tmp(26263) := x"1186";
    tmp(26264) := x"19e8";
    tmp(26265) := x"2aab";
    tmp(26266) := x"53d0";
    tmp(26267) := x"6c93";
    tmp(26268) := x"84f5";
    tmp(26269) := x"a5b7";
    tmp(26270) := x"cf1b";
    tmp(26271) := x"efde";
    tmp(26272) := x"fffd";
    tmp(26273) := x"efd9";
    tmp(26274) := x"ced4";
    tmp(26275) := x"be31";
    tmp(26276) := x"952c";
    tmp(26277) := x"6be7";
    tmp(26278) := x"3a83";
    tmp(26279) := x"21a1";
    tmp(26280) := x"1120";
    tmp(26281) := x"08e0";
    tmp(26282) := x"10e0";
    tmp(26283) := x"1121";
    tmp(26284) := x"29c2";
    tmp(26285) := x"4263";
    tmp(26286) := x"5ae5";
    tmp(26287) := x"7367";
    tmp(26288) := x"83c9";
    tmp(26289) := x"946d";
    tmp(26290) := x"a4f2";
    tmp(26291) := x"9cd3";
    tmp(26292) := x"8c72";
    tmp(26293) := x"740f";
    tmp(26294) := x"634b";
    tmp(26295) := x"4a87";
    tmp(26296) := x"3a04";
    tmp(26297) := x"2982";
    tmp(26298) := x"1921";
    tmp(26299) := x"1921";
    tmp(26300) := x"1101";
    tmp(26301) := x"1921";
    tmp(26302) := x"2181";
    tmp(26303) := x"31e2";
    tmp(26304) := x"4263";
    tmp(26305) := x"5ac4";
    tmp(26306) := x"6b46";
    tmp(26307) := x"7bc7";
    tmp(26308) := x"9c89";
    tmp(26309) := x"b4eb";
    tmp(26310) := x"cd8e";
    tmp(26311) := x"ddee";
    tmp(26312) := x"ee50";
    tmp(26313) := x"e630";
    tmp(26314) := x"d5ef";
    tmp(26315) := x"cd8e";
    tmp(26316) := x"bced";
    tmp(26317) := x"a46b";
    tmp(26318) := x"93ea";
    tmp(26319) := x"83a9";
    tmp(26320) := x"7b88";
    tmp(26321) := x"6b27";
    tmp(26322) := x"6306";
    tmp(26323) := x"5ac6";
    tmp(26324) := x"5285";
    tmp(26325) := x"4a85";
    tmp(26326) := x"4a65";
    tmp(26327) := x"52a5";
    tmp(26328) := x"62e6";
    tmp(26329) := x"7348";
    tmp(26330) := x"8bca";
    tmp(26331) := x"944b";
    tmp(26332) := x"a48d";
    tmp(26333) := x"b52f";
    tmp(26334) := x"bd31";
    tmp(26335) := x"cd92";
    tmp(26336) := x"c572";
    tmp(26337) := x"bd31";
    tmp(26338) := x"acd2";
    tmp(26339) := x"b4d3";
    tmp(26340) := x"b4f5";
    tmp(26341) := x"bcf4";
    tmp(26342) := x"c576";
    tmp(26343) := x"c597";
    tmp(26344) := x"c576";
    tmp(26345) := x"c577";
    tmp(26346) := x"c577";
    tmp(26347) := x"cd78";
    tmp(26348) := x"cd78";
    tmp(26349) := x"cd77";
    tmp(26350) := x"c557";
    tmp(26351) := x"c537";
    tmp(26352) := x"bcd6";
    tmp(26353) := x"bcf6";
    tmp(26354) := x"b4b5";
    tmp(26355) := x"b496";
    tmp(26356) := x"ac75";
    tmp(26357) := x"f800";
    tmp(26358) := x"f800";
    tmp(26359) := x"f800";
    tmp(26360) := x"f800";
    tmp(26361) := x"f800";
    tmp(26362) := x"f800";
    tmp(26363) := x"f800";
    tmp(26364) := x"f800";
    tmp(26365) := x"f800";
    tmp(26366) := x"f800";
    tmp(26367) := x"f800";
    tmp(26368) := x"f800";
    tmp(26369) := x"f800";
    tmp(26370) := x"f800";
    tmp(26371) := x"f800";
    tmp(26372) := x"f800";
    tmp(26373) := x"f800";
    tmp(26374) := x"f800";
    tmp(26375) := x"f800";
    tmp(26376) := x"f800";
    tmp(26377) := x"f800";
    tmp(26378) := x"f800";
    tmp(26379) := x"f800";
    tmp(26380) := x"f800";
    tmp(26381) := x"f800";
    tmp(26382) := x"f800";
    tmp(26383) := x"f800";
    tmp(26384) := x"f800";
    tmp(26385) := x"f800";
    tmp(26386) := x"f800";
    tmp(26387) := x"f800";
    tmp(26388) := x"f800";
    tmp(26389) := x"f800";
    tmp(26390) := x"f800";
    tmp(26391) := x"f800";
    tmp(26392) := x"f800";
    tmp(26393) := x"f800";
    tmp(26394) := x"f800";
    tmp(26395) := x"f800";
    tmp(26396) := x"f800";
    tmp(26397) := x"0840";
    tmp(26398) := x"0840";
    tmp(26399) := x"0840";
    tmp(26400) := x"0020";
    tmp(26401) := x"18c1";
    tmp(26402) := x"10a1";
    tmp(26403) := x"18c1";
    tmp(26404) := x"18e1";
    tmp(26405) := x"18c1";
    tmp(26406) := x"10a1";
    tmp(26407) := x"18a1";
    tmp(26408) := x"20c1";
    tmp(26409) := x"18a1";
    tmp(26410) := x"28c1";
    tmp(26411) := x"49a1";
    tmp(26412) := x"8b63";
    tmp(26413) := x"c4c4";
    tmp(26414) := x"b4a4";
    tmp(26415) := x"7343";
    tmp(26416) := x"4a23";
    tmp(26417) := x"2962";
    tmp(26418) := x"1942";
    tmp(26419) := x"1943";
    tmp(26420) := x"1143";
    tmp(26421) := x"1143";
    tmp(26422) := x"1143";
    tmp(26423) := x"1123";
    tmp(26424) := x"1943";
    tmp(26425) := x"1984";
    tmp(26426) := x"1185";
    tmp(26427) := x"1185";
    tmp(26428) := x"10e3";
    tmp(26429) := x"0861";
    tmp(26430) := x"0904";
    tmp(26431) := x"0924";
    tmp(26432) := x"08e4";
    tmp(26433) := x"08a3";
    tmp(26434) := x"08a3";
    tmp(26435) := x"08e4";
    tmp(26436) := x"08e4";
    tmp(26437) := x"08e4";
    tmp(26438) := x"0905";
    tmp(26439) := x"0905";
    tmp(26440) := x"0905";
    tmp(26441) := x"0904";
    tmp(26442) := x"08a3";
    tmp(26443) := x"08a3";
    tmp(26444) := x"0904";
    tmp(26445) := x"0926";
    tmp(26446) := x"0946";
    tmp(26447) := x"0967";
    tmp(26448) := x"1167";
    tmp(26449) := x"1166";
    tmp(26450) := x"19a6";
    tmp(26451) := x"2163";
    tmp(26452) := x"2921";
    tmp(26453) := x"3100";
    tmp(26454) := x"2921";
    tmp(26455) := x"1102";
    tmp(26456) := x"10e2";
    tmp(26457) := x"08e3";
    tmp(26458) := x"08c3";
    tmp(26459) := x"08c3";
    tmp(26460) := x"08c3";
    tmp(26461) := x"0061";
    tmp(26462) := x"0881";
    tmp(26463) := x"18e1";
    tmp(26464) := x"2920";
    tmp(26465) := x"3960";
    tmp(26466) := x"59e0";
    tmp(26467) := x"7240";
    tmp(26468) := x"8a80";
    tmp(26469) := x"a2e0";
    tmp(26470) := x"b2e0";
    tmp(26471) := x"a2c0";
    tmp(26472) := x"7a80";
    tmp(26473) := x"3181";
    tmp(26474) := x"1122";
    tmp(26475) := x"0903";
    tmp(26476) := x"0924";
    tmp(26477) := x"0904";
    tmp(26478) := x"0924";
    tmp(26479) := x"1145";
    tmp(26480) := x"1165";
    tmp(26481) := x"1144";
    tmp(26482) := x"0924";
    tmp(26483) := x"1144";
    tmp(26484) := x"1165";
    tmp(26485) := x"1164";
    tmp(26486) := x"1164";
    tmp(26487) := x"1144";
    tmp(26488) := x"1123";
    tmp(26489) := x"1123";
    tmp(26490) := x"0924";
    tmp(26491) := x"0944";
    tmp(26492) := x"0965";
    tmp(26493) := x"11a7";
    tmp(26494) := x"09c7";
    tmp(26495) := x"11c7";
    tmp(26496) := x"11c7";
    tmp(26497) := x"1228";
    tmp(26498) := x"1a8a";
    tmp(26499) := x"1208";
    tmp(26500) := x"1166";
    tmp(26501) := x"11a8";
    tmp(26502) := x"330e";
    tmp(26503) := x"6452";
    tmp(26504) := x"95f8";
    tmp(26505) := x"be7a";
    tmp(26506) := x"e75d";
    tmp(26507) := x"ffff";
    tmp(26508) := x"ffff";
    tmp(26509) := x"ffff";
    tmp(26510) := x"ffff";
    tmp(26511) := x"fffe";
    tmp(26512) := x"effb";
    tmp(26513) := x"d736";
    tmp(26514) := x"be72";
    tmp(26515) := x"a5ae";
    tmp(26516) := x"84aa";
    tmp(26517) := x"5b65";
    tmp(26518) := x"2a22";
    tmp(26519) := x"1961";
    tmp(26520) := x"1100";
    tmp(26521) := x"1100";
    tmp(26522) := x"10e0";
    tmp(26523) := x"1100";
    tmp(26524) := x"1961";
    tmp(26525) := x"3202";
    tmp(26526) := x"4264";
    tmp(26527) := x"5b06";
    tmp(26528) := x"7388";
    tmp(26529) := x"8c2c";
    tmp(26530) := x"9cd0";
    tmp(26531) := x"a534";
    tmp(26532) := x"94d3";
    tmp(26533) := x"8450";
    tmp(26534) := x"73cd";
    tmp(26535) := x"5b09";
    tmp(26536) := x"4a86";
    tmp(26537) := x"31e3";
    tmp(26538) := x"2162";
    tmp(26539) := x"1921";
    tmp(26540) := x"1121";
    tmp(26541) := x"1101";
    tmp(26542) := x"1921";
    tmp(26543) := x"2161";
    tmp(26544) := x"29c2";
    tmp(26545) := x"4243";
    tmp(26546) := x"52c4";
    tmp(26547) := x"6325";
    tmp(26548) := x"83e7";
    tmp(26549) := x"9429";
    tmp(26550) := x"acab";
    tmp(26551) := x"cdad";
    tmp(26552) := x"ddef";
    tmp(26553) := x"e630";
    tmp(26554) := x"e630";
    tmp(26555) := x"d5cf";
    tmp(26556) := x"c56e";
    tmp(26557) := x"bd0d";
    tmp(26558) := x"a48b";
    tmp(26559) := x"93ea";
    tmp(26560) := x"8ba9";
    tmp(26561) := x"7b88";
    tmp(26562) := x"7327";
    tmp(26563) := x"62e7";
    tmp(26564) := x"5ac6";
    tmp(26565) := x"5285";
    tmp(26566) := x"4a65";
    tmp(26567) := x"5285";
    tmp(26568) := x"5285";
    tmp(26569) := x"62e7";
    tmp(26570) := x"7348";
    tmp(26571) := x"7bca";
    tmp(26572) := x"8c0b";
    tmp(26573) := x"9c4c";
    tmp(26574) := x"a48d";
    tmp(26575) := x"b4f0";
    tmp(26576) := x"b4f0";
    tmp(26577) := x"a490";
    tmp(26578) := x"a470";
    tmp(26579) := x"acb2";
    tmp(26580) := x"b4d3";
    tmp(26581) := x"bd14";
    tmp(26582) := x"c575";
    tmp(26583) := x"c576";
    tmp(26584) := x"c576";
    tmp(26585) := x"cd97";
    tmp(26586) := x"cd98";
    tmp(26587) := x"cd97";
    tmp(26588) := x"c577";
    tmp(26589) := x"c557";
    tmp(26590) := x"c517";
    tmp(26591) := x"bcf7";
    tmp(26592) := x"b4b6";
    tmp(26593) := x"b4b5";
    tmp(26594) := x"ac95";
    tmp(26595) := x"ac55";
    tmp(26596) := x"a475";
    tmp(26597) := x"f800";
    tmp(26598) := x"f800";
    tmp(26599) := x"f800";
    tmp(26600) := x"f800";
    tmp(26601) := x"f800";
    tmp(26602) := x"f800";
    tmp(26603) := x"f800";
    tmp(26604) := x"f800";
    tmp(26605) := x"f800";
    tmp(26606) := x"f800";
    tmp(26607) := x"f800";
    tmp(26608) := x"f800";
    tmp(26609) := x"f800";
    tmp(26610) := x"f800";
    tmp(26611) := x"f800";
    tmp(26612) := x"f800";
    tmp(26613) := x"f800";
    tmp(26614) := x"f800";
    tmp(26615) := x"f800";
    tmp(26616) := x"f800";
    tmp(26617) := x"f800";
    tmp(26618) := x"f800";
    tmp(26619) := x"f800";
    tmp(26620) := x"f800";
    tmp(26621) := x"f800";
    tmp(26622) := x"f800";
    tmp(26623) := x"f800";
    tmp(26624) := x"f800";
    tmp(26625) := x"f800";
    tmp(26626) := x"f800";
    tmp(26627) := x"f800";
    tmp(26628) := x"f800";
    tmp(26629) := x"f800";
    tmp(26630) := x"f800";
    tmp(26631) := x"f800";
    tmp(26632) := x"f800";
    tmp(26633) := x"f800";
    tmp(26634) := x"f800";
    tmp(26635) := x"f800";
    tmp(26636) := x"f800";
    tmp(26637) := x"0860";
    tmp(26638) := x"0840";
    tmp(26639) := x"0840";
    tmp(26640) := x"0020";
    tmp(26641) := x"1924";
    tmp(26642) := x"1944";
    tmp(26643) := x"1923";
    tmp(26644) := x"1924";
    tmp(26645) := x"2144";
    tmp(26646) := x"2943";
    tmp(26647) := x"3183";
    tmp(26648) := x"3142";
    tmp(26649) := x"20e1";
    tmp(26650) := x"20e1";
    tmp(26651) := x"2902";
    tmp(26652) := x"3961";
    tmp(26653) := x"6262";
    tmp(26654) := x"8343";
    tmp(26655) := x"bd26";
    tmp(26656) := x"6367";
    tmp(26657) := x"1125";
    tmp(26658) := x"0926";
    tmp(26659) := x"0925";
    tmp(26660) := x"0925";
    tmp(26661) := x"0905";
    tmp(26662) := x"0905";
    tmp(26663) := x"08e5";
    tmp(26664) := x"0905";
    tmp(26665) := x"0905";
    tmp(26666) := x"0905";
    tmp(26667) := x"0905";
    tmp(26668) := x"08a3";
    tmp(26669) := x"0041";
    tmp(26670) := x"0041";
    tmp(26671) := x"08a3";
    tmp(26672) := x"08a3";
    tmp(26673) := x"08a3";
    tmp(26674) := x"08c4";
    tmp(26675) := x"08e4";
    tmp(26676) := x"08e5";
    tmp(26677) := x"08e5";
    tmp(26678) := x"08e4";
    tmp(26679) := x"08e4";
    tmp(26680) := x"0905";
    tmp(26681) := x"08c3";
    tmp(26682) := x"0041";
    tmp(26683) := x"0041";
    tmp(26684) := x"0062";
    tmp(26685) := x"08e4";
    tmp(26686) := x"0925";
    tmp(26687) := x"0926";
    tmp(26688) := x"0926";
    tmp(26689) := x"1166";
    tmp(26690) := x"1187";
    tmp(26691) := x"19c8";
    tmp(26692) := x"10c3";
    tmp(26693) := x"1061";
    tmp(26694) := x"10a1";
    tmp(26695) := x"08a3";
    tmp(26696) := x"08c3";
    tmp(26697) := x"08c3";
    tmp(26698) := x"08a3";
    tmp(26699) := x"00a2";
    tmp(26700) := x"0061";
    tmp(26701) := x"0041";
    tmp(26702) := x"08a2";
    tmp(26703) := x"08c2";
    tmp(26704) := x"1901";
    tmp(26705) := x"3161";
    tmp(26706) := x"49e0";
    tmp(26707) := x"5a00";
    tmp(26708) := x"6a40";
    tmp(26709) := x"7260";
    tmp(26710) := x"7a80";
    tmp(26711) := x"5a20";
    tmp(26712) := x"2981";
    tmp(26713) := x"1102";
    tmp(26714) := x"0903";
    tmp(26715) := x"0904";
    tmp(26716) := x"0924";
    tmp(26717) := x"0925";
    tmp(26718) := x"0966";
    tmp(26719) := x"11c7";
    tmp(26720) := x"11a7";
    tmp(26721) := x"0945";
    tmp(26722) := x"0966";
    tmp(26723) := x"1186";
    tmp(26724) := x"1186";
    tmp(26725) := x"1186";
    tmp(26726) := x"0965";
    tmp(26727) := x"0945";
    tmp(26728) := x"0904";
    tmp(26729) := x"0924";
    tmp(26730) := x"0965";
    tmp(26731) := x"1186";
    tmp(26732) := x"11c7";
    tmp(26733) := x"11a6";
    tmp(26734) := x"11e7";
    tmp(26735) := x"11e7";
    tmp(26736) := x"11c7";
    tmp(26737) := x"1186";
    tmp(26738) := x"1166";
    tmp(26739) := x"2a4a";
    tmp(26740) := x"6c53";
    tmp(26741) := x"b639";
    tmp(26742) := x"d71c";
    tmp(26743) := x"ef9e";
    tmp(26744) := x"ffff";
    tmp(26745) := x"ffff";
    tmp(26746) := x"ffff";
    tmp(26747) := x"ffff";
    tmp(26748) := x"ffff";
    tmp(26749) := x"ffff";
    tmp(26750) := x"ffff";
    tmp(26751) := x"f7fd";
    tmp(26752) := x"e799";
    tmp(26753) := x"cef5";
    tmp(26754) := x"adf0";
    tmp(26755) := x"8d2b";
    tmp(26756) := x"63c6";
    tmp(26757) := x"42e3";
    tmp(26758) := x"21c1";
    tmp(26759) := x"1120";
    tmp(26760) := x"1100";
    tmp(26761) := x"1100";
    tmp(26762) := x"1100";
    tmp(26763) := x"1100";
    tmp(26764) := x"1120";
    tmp(26765) := x"2181";
    tmp(26766) := x"3202";
    tmp(26767) := x"4a84";
    tmp(26768) := x"6326";
    tmp(26769) := x"7bca";
    tmp(26770) := x"948e";
    tmp(26771) := x"9cf1";
    tmp(26772) := x"94f3";
    tmp(26773) := x"94d2";
    tmp(26774) := x"73ee";
    tmp(26775) := x"6b6b";
    tmp(26776) := x"52a7";
    tmp(26777) := x"4a65";
    tmp(26778) := x"31e3";
    tmp(26779) := x"2162";
    tmp(26780) := x"1921";
    tmp(26781) := x"1101";
    tmp(26782) := x"1101";
    tmp(26783) := x"1921";
    tmp(26784) := x"2161";
    tmp(26785) := x"29a2";
    tmp(26786) := x"3a22";
    tmp(26787) := x"52a4";
    tmp(26788) := x"6b25";
    tmp(26789) := x"7b87";
    tmp(26790) := x"9429";
    tmp(26791) := x"b4cb";
    tmp(26792) := x"c56d";
    tmp(26793) := x"ddef";
    tmp(26794) := x"e630";
    tmp(26795) := x"de10";
    tmp(26796) := x"cdaf";
    tmp(26797) := x"c54e";
    tmp(26798) := x"b4cd";
    tmp(26799) := x"a48b";
    tmp(26800) := x"940a";
    tmp(26801) := x"83c9";
    tmp(26802) := x"7b89";
    tmp(26803) := x"7348";
    tmp(26804) := x"6307";
    tmp(26805) := x"5ac6";
    tmp(26806) := x"5285";
    tmp(26807) := x"5285";
    tmp(26808) := x"52a5";
    tmp(26809) := x"5ac6";
    tmp(26810) := x"6307";
    tmp(26811) := x"6b28";
    tmp(26812) := x"7369";
    tmp(26813) := x"8bcb";
    tmp(26814) := x"940c";
    tmp(26815) := x"9c4d";
    tmp(26816) := x"a44e";
    tmp(26817) := x"93ee";
    tmp(26818) := x"9c4f";
    tmp(26819) := x"a451";
    tmp(26820) := x"ac92";
    tmp(26821) := x"bcf3";
    tmp(26822) := x"bd35";
    tmp(26823) := x"c576";
    tmp(26824) := x"c577";
    tmp(26825) := x"c557";
    tmp(26826) := x"cd98";
    tmp(26827) := x"cdb7";
    tmp(26828) := x"c577";
    tmp(26829) := x"c537";
    tmp(26830) := x"bcf7";
    tmp(26831) := x"bcd6";
    tmp(26832) := x"b4b6";
    tmp(26833) := x"acb6";
    tmp(26834) := x"a495";
    tmp(26835) := x"ac96";
    tmp(26836) := x"a475";
    tmp(26837) := x"f800";
    tmp(26838) := x"f800";
    tmp(26839) := x"f800";
    tmp(26840) := x"f800";
    tmp(26841) := x"f800";
    tmp(26842) := x"f800";
    tmp(26843) := x"f800";
    tmp(26844) := x"f800";
    tmp(26845) := x"f800";
    tmp(26846) := x"f800";
    tmp(26847) := x"f800";
    tmp(26848) := x"f800";
    tmp(26849) := x"f800";
    tmp(26850) := x"f800";
    tmp(26851) := x"f800";
    tmp(26852) := x"f800";
    tmp(26853) := x"f800";
    tmp(26854) := x"f800";
    tmp(26855) := x"f800";
    tmp(26856) := x"f800";
    tmp(26857) := x"f800";
    tmp(26858) := x"f800";
    tmp(26859) := x"f800";
    tmp(26860) := x"f800";
    tmp(26861) := x"f800";
    tmp(26862) := x"f800";
    tmp(26863) := x"f800";
    tmp(26864) := x"f800";
    tmp(26865) := x"f800";
    tmp(26866) := x"f800";
    tmp(26867) := x"f800";
    tmp(26868) := x"f800";
    tmp(26869) := x"f800";
    tmp(26870) := x"f800";
    tmp(26871) := x"f800";
    tmp(26872) := x"f800";
    tmp(26873) := x"f800";
    tmp(26874) := x"f800";
    tmp(26875) := x"f800";
    tmp(26876) := x"f800";
    tmp(26877) := x"0861";
    tmp(26878) := x"0840";
    tmp(26879) := x"0840";
    tmp(26880) := x"0020";
    tmp(26881) := x"1904";
    tmp(26882) := x"1924";
    tmp(26883) := x"10a3";
    tmp(26884) := x"10a3";
    tmp(26885) := x"10a2";
    tmp(26886) := x"0861";
    tmp(26887) := x"0861";
    tmp(26888) := x"1081";
    tmp(26889) := x"20e2";
    tmp(26890) := x"3984";
    tmp(26891) := x"5225";
    tmp(26892) := x"62a7";
    tmp(26893) := x"6287";
    tmp(26894) := x"6ae8";
    tmp(26895) := x"39c5";
    tmp(26896) := x"10e3";
    tmp(26897) := x"0883";
    tmp(26898) := x"08a4";
    tmp(26899) := x"08e4";
    tmp(26900) := x"08a3";
    tmp(26901) := x"0062";
    tmp(26902) := x"0041";
    tmp(26903) := x"0041";
    tmp(26904) := x"0082";
    tmp(26905) := x"00a4";
    tmp(26906) := x"00a4";
    tmp(26907) := x"00a4";
    tmp(26908) := x"08c4";
    tmp(26909) := x"08a4";
    tmp(26910) := x"0882";
    tmp(26911) := x"00a3";
    tmp(26912) := x"08c4";
    tmp(26913) := x"08e4";
    tmp(26914) := x"08e5";
    tmp(26915) := x"08c4";
    tmp(26916) := x"08c4";
    tmp(26917) := x"0905";
    tmp(26918) := x"0925";
    tmp(26919) := x"0905";
    tmp(26920) := x"0905";
    tmp(26921) := x"08a3";
    tmp(26922) := x"08a3";
    tmp(26923) := x"0882";
    tmp(26924) := x"08a3";
    tmp(26925) := x"08e4";
    tmp(26926) := x"08c4";
    tmp(26927) := x"08e4";
    tmp(26928) := x"08e4";
    tmp(26929) := x"08c4";
    tmp(26930) := x"08a3";
    tmp(26931) := x"08c4";
    tmp(26932) := x"08a2";
    tmp(26933) := x"0861";
    tmp(26934) := x"10e3";
    tmp(26935) := x"08e3";
    tmp(26936) := x"00a2";
    tmp(26937) := x"0082";
    tmp(26938) := x"0061";
    tmp(26939) := x"0041";
    tmp(26940) := x"0082";
    tmp(26941) := x"0904";
    tmp(26942) := x"0905";
    tmp(26943) := x"08c3";
    tmp(26944) := x"08e2";
    tmp(26945) := x"1942";
    tmp(26946) := x"2142";
    tmp(26947) := x"2161";
    tmp(26948) := x"3160";
    tmp(26949) := x"41a0";
    tmp(26950) := x"49e0";
    tmp(26951) := x"2981";
    tmp(26952) := x"1142";
    tmp(26953) := x"0903";
    tmp(26954) := x"0904";
    tmp(26955) := x"0924";
    tmp(26956) := x"0966";
    tmp(26957) := x"11a7";
    tmp(26958) := x"1187";
    tmp(26959) := x"1187";
    tmp(26960) := x"1166";
    tmp(26961) := x"0966";
    tmp(26962) := x"0946";
    tmp(26963) := x"0946";
    tmp(26964) := x"0965";
    tmp(26965) := x"0945";
    tmp(26966) := x"0945";
    tmp(26967) := x"0925";
    tmp(26968) := x"0965";
    tmp(26969) := x"0986";
    tmp(26970) := x"11c7";
    tmp(26971) := x"1208";
    tmp(26972) := x"11e8";
    tmp(26973) := x"11c7";
    tmp(26974) := x"1186";
    tmp(26975) := x"1165";
    tmp(26976) := x"1124";
    tmp(26977) := x"2187";
    tmp(26978) := x"6c32";
    tmp(26979) := x"cedb";
    tmp(26980) := x"f7bf";
    tmp(26981) := x"ffff";
    tmp(26982) := x"ffff";
    tmp(26983) := x"ffff";
    tmp(26984) := x"ffff";
    tmp(26985) := x"ffff";
    tmp(26986) := x"ffff";
    tmp(26987) := x"ffff";
    tmp(26988) := x"ffff";
    tmp(26989) := x"ffff";
    tmp(26990) := x"ffff";
    tmp(26991) := x"f7fb";
    tmp(26992) := x"df97";
    tmp(26993) := x"be52";
    tmp(26994) := x"956d";
    tmp(26995) := x"7428";
    tmp(26996) := x"4b24";
    tmp(26997) := x"3242";
    tmp(26998) := x"19a1";
    tmp(26999) := x"1120";
    tmp(27000) := x"1120";
    tmp(27001) := x"1100";
    tmp(27002) := x"1100";
    tmp(27003) := x"1100";
    tmp(27004) := x"1100";
    tmp(27005) := x"1121";
    tmp(27006) := x"21a1";
    tmp(27007) := x"3a23";
    tmp(27008) := x"52c5";
    tmp(27009) := x"6b88";
    tmp(27010) := x"844c";
    tmp(27011) := x"8c8f";
    tmp(27012) := x"9cf2";
    tmp(27013) := x"94f2";
    tmp(27014) := x"8c8f";
    tmp(27015) := x"7bec";
    tmp(27016) := x"6349";
    tmp(27017) := x"52a6";
    tmp(27018) := x"4224";
    tmp(27019) := x"29a2";
    tmp(27020) := x"2161";
    tmp(27021) := x"1921";
    tmp(27022) := x"1101";
    tmp(27023) := x"1101";
    tmp(27024) := x"1921";
    tmp(27025) := x"2161";
    tmp(27026) := x"29a1";
    tmp(27027) := x"4223";
    tmp(27028) := x"52a4";
    tmp(27029) := x"6b26";
    tmp(27030) := x"7b87";
    tmp(27031) := x"9449";
    tmp(27032) := x"accb";
    tmp(27033) := x"c56d";
    tmp(27034) := x"d5ae";
    tmp(27035) := x"d5ef";
    tmp(27036) := x"cdae";
    tmp(27037) := x"cd6e";
    tmp(27038) := x"c54e";
    tmp(27039) := x"b4cc";
    tmp(27040) := x"a46c";
    tmp(27041) := x"940b";
    tmp(27042) := x"8c0a";
    tmp(27043) := x"7b89";
    tmp(27044) := x"6b48";
    tmp(27045) := x"6307";
    tmp(27046) := x"5ae6";
    tmp(27047) := x"5285";
    tmp(27048) := x"5285";
    tmp(27049) := x"52a6";
    tmp(27050) := x"5ac7";
    tmp(27051) := x"62e7";
    tmp(27052) := x"6b28";
    tmp(27053) := x"736a";
    tmp(27054) := x"7b6b";
    tmp(27055) := x"838b";
    tmp(27056) := x"838c";
    tmp(27057) := x"8bad";
    tmp(27058) := x"93ee";
    tmp(27059) := x"9410";
    tmp(27060) := x"ac72";
    tmp(27061) := x"b4f3";
    tmp(27062) := x"c576";
    tmp(27063) := x"bd37";
    tmp(27064) := x"c578";
    tmp(27065) := x"c578";
    tmp(27066) := x"cd99";
    tmp(27067) := x"c577";
    tmp(27068) := x"c557";
    tmp(27069) := x"bcf6";
    tmp(27070) := x"bcf8";
    tmp(27071) := x"b4f8";
    tmp(27072) := x"b4b7";
    tmp(27073) := x"ac95";
    tmp(27074) := x"ac75";
    tmp(27075) := x"ac96";
    tmp(27076) := x"a475";
    tmp(27077) := x"f800";
    tmp(27078) := x"f800";
    tmp(27079) := x"f800";
    tmp(27080) := x"f800";
    tmp(27081) := x"f800";
    tmp(27082) := x"f800";
    tmp(27083) := x"f800";
    tmp(27084) := x"f800";
    tmp(27085) := x"f800";
    tmp(27086) := x"f800";
    tmp(27087) := x"f800";
    tmp(27088) := x"f800";
    tmp(27089) := x"f800";
    tmp(27090) := x"f800";
    tmp(27091) := x"f800";
    tmp(27092) := x"f800";
    tmp(27093) := x"f800";
    tmp(27094) := x"f800";
    tmp(27095) := x"f800";
    tmp(27096) := x"f800";
    tmp(27097) := x"f800";
    tmp(27098) := x"f800";
    tmp(27099) := x"f800";
    tmp(27100) := x"f800";
    tmp(27101) := x"f800";
    tmp(27102) := x"f800";
    tmp(27103) := x"f800";
    tmp(27104) := x"f800";
    tmp(27105) := x"f800";
    tmp(27106) := x"f800";
    tmp(27107) := x"f800";
    tmp(27108) := x"f800";
    tmp(27109) := x"f800";
    tmp(27110) := x"f800";
    tmp(27111) := x"f800";
    tmp(27112) := x"f800";
    tmp(27113) := x"f800";
    tmp(27114) := x"f800";
    tmp(27115) := x"f800";
    tmp(27116) := x"f800";
    tmp(27117) := x"0840";
    tmp(27118) := x"0860";
    tmp(27119) := x"0840";
    tmp(27120) := x"0000";
    tmp(27121) := x"0884";
    tmp(27122) := x"0864";
    tmp(27123) := x"0063";
    tmp(27124) := x"0063";
    tmp(27125) := x"0043";
    tmp(27126) := x"0043";
    tmp(27127) := x"0042";
    tmp(27128) := x"0862";
    tmp(27129) := x"10a3";
    tmp(27130) := x"1904";
    tmp(27131) := x"2945";
    tmp(27132) := x"31a7";
    tmp(27133) := x"31a7";
    tmp(27134) := x"3186";
    tmp(27135) := x"10a3";
    tmp(27136) := x"08a3";
    tmp(27137) := x"08a3";
    tmp(27138) := x"0062";
    tmp(27139) := x"0021";
    tmp(27140) := x"0020";
    tmp(27141) := x"0021";
    tmp(27142) := x"0041";
    tmp(27143) := x"0062";
    tmp(27144) := x"0082";
    tmp(27145) := x"00a3";
    tmp(27146) := x"00a4";
    tmp(27147) := x"00c4";
    tmp(27148) := x"00a4";
    tmp(27149) := x"00a4";
    tmp(27150) := x"08c4";
    tmp(27151) := x"08e5";
    tmp(27152) := x"08c4";
    tmp(27153) := x"08c4";
    tmp(27154) := x"08c4";
    tmp(27155) := x"08a3";
    tmp(27156) := x"08c4";
    tmp(27157) := x"08e4";
    tmp(27158) := x"08c4";
    tmp(27159) := x"08c4";
    tmp(27160) := x"08c4";
    tmp(27161) := x"0062";
    tmp(27162) := x"0882";
    tmp(27163) := x"0882";
    tmp(27164) := x"08c4";
    tmp(27165) := x"08e5";
    tmp(27166) := x"0905";
    tmp(27167) := x"08e4";
    tmp(27168) := x"0925";
    tmp(27169) := x"08e4";
    tmp(27170) := x"08a3";
    tmp(27171) := x"08c3";
    tmp(27172) := x"0882";
    tmp(27173) := x"0861";
    tmp(27174) := x"1104";
    tmp(27175) := x"1186";
    tmp(27176) := x"08c3";
    tmp(27177) := x"0041";
    tmp(27178) := x"0061";
    tmp(27179) := x"08c3";
    tmp(27180) := x"0946";
    tmp(27181) := x"0926";
    tmp(27182) := x"0905";
    tmp(27183) := x"0904";
    tmp(27184) := x"0904";
    tmp(27185) := x"0905";
    tmp(27186) := x"08e4";
    tmp(27187) := x"08e2";
    tmp(27188) := x"1901";
    tmp(27189) := x"2141";
    tmp(27190) := x"1981";
    tmp(27191) := x"1163";
    tmp(27192) := x"0924";
    tmp(27193) := x"0924";
    tmp(27194) := x"0945";
    tmp(27195) := x"11a7";
    tmp(27196) := x"11e8";
    tmp(27197) := x"11a7";
    tmp(27198) := x"0966";
    tmp(27199) := x"0945";
    tmp(27200) := x"0924";
    tmp(27201) := x"0904";
    tmp(27202) := x"0904";
    tmp(27203) := x"0904";
    tmp(27204) := x"0904";
    tmp(27205) := x"0924";
    tmp(27206) := x"0965";
    tmp(27207) := x"0966";
    tmp(27208) := x"1186";
    tmp(27209) := x"11a7";
    tmp(27210) := x"11c8";
    tmp(27211) := x"19e8";
    tmp(27212) := x"11a6";
    tmp(27213) := x"1145";
    tmp(27214) := x"1146";
    tmp(27215) := x"29e9";
    tmp(27216) := x"7433";
    tmp(27217) := x"d6fd";
    tmp(27218) := x"ffdf";
    tmp(27219) := x"ffff";
    tmp(27220) := x"ffff";
    tmp(27221) := x"ffff";
    tmp(27222) := x"ffff";
    tmp(27223) := x"ffff";
    tmp(27224) := x"ffff";
    tmp(27225) := x"ffff";
    tmp(27226) := x"ffff";
    tmp(27227) := x"ffff";
    tmp(27228) := x"ffff";
    tmp(27229) := x"ffff";
    tmp(27230) := x"fffe";
    tmp(27231) := x"effb";
    tmp(27232) := x"cf35";
    tmp(27233) := x"adef";
    tmp(27234) := x"7cca";
    tmp(27235) := x"5365";
    tmp(27236) := x"3a82";
    tmp(27237) := x"21c1";
    tmp(27238) := x"1961";
    tmp(27239) := x"1141";
    tmp(27240) := x"1141";
    tmp(27241) := x"1121";
    tmp(27242) := x"1120";
    tmp(27243) := x"1120";
    tmp(27244) := x"1100";
    tmp(27245) := x"1100";
    tmp(27246) := x"1921";
    tmp(27247) := x"29c2";
    tmp(27248) := x"4264";
    tmp(27249) := x"5b47";
    tmp(27250) := x"73aa";
    tmp(27251) := x"842c";
    tmp(27252) := x"8caf";
    tmp(27253) := x"94d0";
    tmp(27254) := x"94f0";
    tmp(27255) := x"8c4e";
    tmp(27256) := x"73aa";
    tmp(27257) := x"6348";
    tmp(27258) := x"4a85";
    tmp(27259) := x"3a04";
    tmp(27260) := x"29a2";
    tmp(27261) := x"2141";
    tmp(27262) := x"1921";
    tmp(27263) := x"1101";
    tmp(27264) := x"1921";
    tmp(27265) := x"1921";
    tmp(27266) := x"2161";
    tmp(27267) := x"31c2";
    tmp(27268) := x"3a02";
    tmp(27269) := x"5284";
    tmp(27270) := x"6305";
    tmp(27271) := x"7387";
    tmp(27272) := x"9409";
    tmp(27273) := x"accb";
    tmp(27274) := x"c52d";
    tmp(27275) := x"cdae";
    tmp(27276) := x"cd8e";
    tmp(27277) := x"c56e";
    tmp(27278) := x"c52e";
    tmp(27279) := x"b4ed";
    tmp(27280) := x"b4cd";
    tmp(27281) := x"a46c";
    tmp(27282) := x"940b";
    tmp(27283) := x"83ca";
    tmp(27284) := x"7ba9";
    tmp(27285) := x"7368";
    tmp(27286) := x"6b07";
    tmp(27287) := x"5ac6";
    tmp(27288) := x"5286";
    tmp(27289) := x"52a6";
    tmp(27290) := x"52a7";
    tmp(27291) := x"5aa7";
    tmp(27292) := x"62c8";
    tmp(27293) := x"6b29";
    tmp(27294) := x"734a";
    tmp(27295) := x"7b6a";
    tmp(27296) := x"7b4a";
    tmp(27297) := x"838c";
    tmp(27298) := x"8bad";
    tmp(27299) := x"93ef";
    tmp(27300) := x"a472";
    tmp(27301) := x"acd2";
    tmp(27302) := x"bd35";
    tmp(27303) := x"bd37";
    tmp(27304) := x"c577";
    tmp(27305) := x"c578";
    tmp(27306) := x"cd99";
    tmp(27307) := x"c578";
    tmp(27308) := x"bd37";
    tmp(27309) := x"b4d6";
    tmp(27310) := x"bcf7";
    tmp(27311) := x"b4f7";
    tmp(27312) := x"b4b6";
    tmp(27313) := x"b476";
    tmp(27314) := x"ac95";
    tmp(27315) := x"ac75";
    tmp(27316) := x"ac76";
    tmp(27317) := x"f800";
    tmp(27318) := x"f800";
    tmp(27319) := x"f800";
    tmp(27320) := x"f800";
    tmp(27321) := x"f800";
    tmp(27322) := x"f800";
    tmp(27323) := x"f800";
    tmp(27324) := x"f800";
    tmp(27325) := x"f800";
    tmp(27326) := x"f800";
    tmp(27327) := x"f800";
    tmp(27328) := x"f800";
    tmp(27329) := x"f800";
    tmp(27330) := x"f800";
    tmp(27331) := x"f800";
    tmp(27332) := x"f800";
    tmp(27333) := x"f800";
    tmp(27334) := x"f800";
    tmp(27335) := x"f800";
    tmp(27336) := x"f800";
    tmp(27337) := x"f800";
    tmp(27338) := x"f800";
    tmp(27339) := x"f800";
    tmp(27340) := x"f800";
    tmp(27341) := x"f800";
    tmp(27342) := x"f800";
    tmp(27343) := x"f800";
    tmp(27344) := x"f800";
    tmp(27345) := x"f800";
    tmp(27346) := x"f800";
    tmp(27347) := x"f800";
    tmp(27348) := x"f800";
    tmp(27349) := x"f800";
    tmp(27350) := x"f800";
    tmp(27351) := x"f800";
    tmp(27352) := x"f800";
    tmp(27353) := x"f800";
    tmp(27354) := x"f800";
    tmp(27355) := x"f800";
    tmp(27356) := x"f800";
    tmp(27357) := x"0840";
    tmp(27358) := x"0840";
    tmp(27359) := x"0860";
    tmp(27360) := x"0000";
    tmp(27361) := x"0044";
    tmp(27362) := x"0044";
    tmp(27363) := x"0044";
    tmp(27364) := x"0044";
    tmp(27365) := x"0044";
    tmp(27366) := x"0044";
    tmp(27367) := x"0044";
    tmp(27368) := x"0043";
    tmp(27369) := x"0043";
    tmp(27370) := x"0043";
    tmp(27371) := x"0043";
    tmp(27372) := x"0843";
    tmp(27373) := x"0843";
    tmp(27374) := x"0842";
    tmp(27375) := x"0020";
    tmp(27376) := x"0021";
    tmp(27377) := x"0041";
    tmp(27378) := x"0041";
    tmp(27379) := x"0021";
    tmp(27380) := x"0041";
    tmp(27381) := x"0062";
    tmp(27382) := x"0083";
    tmp(27383) := x"00a3";
    tmp(27384) := x"00a4";
    tmp(27385) := x"00a4";
    tmp(27386) := x"00a4";
    tmp(27387) := x"00a3";
    tmp(27388) := x"00c4";
    tmp(27389) := x"08e5";
    tmp(27390) := x"08c4";
    tmp(27391) := x"08c4";
    tmp(27392) := x"00a3";
    tmp(27393) := x"08a3";
    tmp(27394) := x"08a3";
    tmp(27395) := x"08c4";
    tmp(27396) := x"08c4";
    tmp(27397) := x"08c4";
    tmp(27398) := x"08c4";
    tmp(27399) := x"08c4";
    tmp(27400) := x"08c4";
    tmp(27401) := x"0883";
    tmp(27402) := x"08a3";
    tmp(27403) := x"08a3";
    tmp(27404) := x"08c4";
    tmp(27405) := x"08c4";
    tmp(27406) := x"08e4";
    tmp(27407) := x"0904";
    tmp(27408) := x"0905";
    tmp(27409) := x"08c3";
    tmp(27410) := x"08c4";
    tmp(27411) := x"08e4";
    tmp(27412) := x"08c3";
    tmp(27413) := x"0882";
    tmp(27414) := x"10e4";
    tmp(27415) := x"1166";
    tmp(27416) := x"1166";
    tmp(27417) := x"0904";
    tmp(27418) := x"0904";
    tmp(27419) := x"0926";
    tmp(27420) := x"0946";
    tmp(27421) := x"0926";
    tmp(27422) := x"0926";
    tmp(27423) := x"0926";
    tmp(27424) := x"0925";
    tmp(27425) := x"0926";
    tmp(27426) := x"0925";
    tmp(27427) := x"0925";
    tmp(27428) := x"1124";
    tmp(27429) := x"1103";
    tmp(27430) := x"1123";
    tmp(27431) := x"1164";
    tmp(27432) := x"1185";
    tmp(27433) := x"1186";
    tmp(27434) := x"1187";
    tmp(27435) := x"0966";
    tmp(27436) := x"0945";
    tmp(27437) := x"0945";
    tmp(27438) := x"0925";
    tmp(27439) := x"0904";
    tmp(27440) := x"0904";
    tmp(27441) := x"0904";
    tmp(27442) := x"0924";
    tmp(27443) := x"0924";
    tmp(27444) := x"0965";
    tmp(27445) := x"11a6";
    tmp(27446) := x"11a7";
    tmp(27447) := x"1146";
    tmp(27448) := x"1145";
    tmp(27449) := x"1946";
    tmp(27450) := x"21a8";
    tmp(27451) := x"2a0a";
    tmp(27452) := x"42cd";
    tmp(27453) := x"7c73";
    tmp(27454) := x"c65c";
    tmp(27455) := x"f7df";
    tmp(27456) := x"ffdf";
    tmp(27457) := x"ffff";
    tmp(27458) := x"ffff";
    tmp(27459) := x"ffff";
    tmp(27460) := x"ffff";
    tmp(27461) := x"ffff";
    tmp(27462) := x"ffff";
    tmp(27463) := x"ffff";
    tmp(27464) := x"ffff";
    tmp(27465) := x"ffff";
    tmp(27466) := x"ffff";
    tmp(27467) := x"ffff";
    tmp(27468) := x"ffff";
    tmp(27469) := x"ffff";
    tmp(27470) := x"f7dc";
    tmp(27471) := x"df57";
    tmp(27472) := x"b631";
    tmp(27473) := x"84ec";
    tmp(27474) := x"5ba7";
    tmp(27475) := x"3aa3";
    tmp(27476) := x"2a01";
    tmp(27477) := x"1961";
    tmp(27478) := x"1140";
    tmp(27479) := x"1981";
    tmp(27480) := x"1961";
    tmp(27481) := x"1121";
    tmp(27482) := x"1121";
    tmp(27483) := x"1121";
    tmp(27484) := x"1101";
    tmp(27485) := x"1101";
    tmp(27486) := x"1101";
    tmp(27487) := x"1961";
    tmp(27488) := x"31e2";
    tmp(27489) := x"4aa4";
    tmp(27490) := x"6b88";
    tmp(27491) := x"7beb";
    tmp(27492) := x"8c6d";
    tmp(27493) := x"8c8e";
    tmp(27494) := x"94ae";
    tmp(27495) := x"9ccf";
    tmp(27496) := x"83eb";
    tmp(27497) := x"738a";
    tmp(27498) := x"5ae7";
    tmp(27499) := x"4a65";
    tmp(27500) := x"39e3";
    tmp(27501) := x"2982";
    tmp(27502) := x"2141";
    tmp(27503) := x"1921";
    tmp(27504) := x"1101";
    tmp(27505) := x"1901";
    tmp(27506) := x"1921";
    tmp(27507) := x"2141";
    tmp(27508) := x"31a2";
    tmp(27509) := x"4222";
    tmp(27510) := x"5284";
    tmp(27511) := x"62e5";
    tmp(27512) := x"7b87";
    tmp(27513) := x"9449";
    tmp(27514) := x"accb";
    tmp(27515) := x"bd4d";
    tmp(27516) := x"cdae";
    tmp(27517) := x"c54d";
    tmp(27518) := x"c52d";
    tmp(27519) := x"bced";
    tmp(27520) := x"b4cd";
    tmp(27521) := x"ac8d";
    tmp(27522) := x"a46c";
    tmp(27523) := x"942b";
    tmp(27524) := x"8c0b";
    tmp(27525) := x"7b89";
    tmp(27526) := x"7b89";
    tmp(27527) := x"6b07";
    tmp(27528) := x"5ac6";
    tmp(27529) := x"5286";
    tmp(27530) := x"5266";
    tmp(27531) := x"5286";
    tmp(27532) := x"5aa7";
    tmp(27533) := x"62c8";
    tmp(27534) := x"6ae8";
    tmp(27535) := x"7329";
    tmp(27536) := x"6b09";
    tmp(27537) := x"7b4a";
    tmp(27538) := x"838d";
    tmp(27539) := x"93ef";
    tmp(27540) := x"9c31";
    tmp(27541) := x"a492";
    tmp(27542) := x"b4f4";
    tmp(27543) := x"c557";
    tmp(27544) := x"bd57";
    tmp(27545) := x"bd78";
    tmp(27546) := x"bd58";
    tmp(27547) := x"bd38";
    tmp(27548) := x"b4d7";
    tmp(27549) := x"acb7";
    tmp(27550) := x"b4d6";
    tmp(27551) := x"b4d6";
    tmp(27552) := x"b496";
    tmp(27553) := x"ac95";
    tmp(27554) := x"a454";
    tmp(27555) := x"a455";
    tmp(27556) := x"a415";
    tmp(27557) := x"f800";
    tmp(27558) := x"f800";
    tmp(27559) := x"f800";
    tmp(27560) := x"f800";
    tmp(27561) := x"f800";
    tmp(27562) := x"f800";
    tmp(27563) := x"f800";
    tmp(27564) := x"f800";
    tmp(27565) := x"f800";
    tmp(27566) := x"f800";
    tmp(27567) := x"f800";
    tmp(27568) := x"f800";
    tmp(27569) := x"f800";
    tmp(27570) := x"f800";
    tmp(27571) := x"f800";
    tmp(27572) := x"f800";
    tmp(27573) := x"f800";
    tmp(27574) := x"f800";
    tmp(27575) := x"f800";
    tmp(27576) := x"f800";
    tmp(27577) := x"f800";
    tmp(27578) := x"f800";
    tmp(27579) := x"f800";
    tmp(27580) := x"f800";
    tmp(27581) := x"f800";
    tmp(27582) := x"f800";
    tmp(27583) := x"f800";
    tmp(27584) := x"f800";
    tmp(27585) := x"f800";
    tmp(27586) := x"f800";
    tmp(27587) := x"f800";
    tmp(27588) := x"f800";
    tmp(27589) := x"f800";
    tmp(27590) := x"f800";
    tmp(27591) := x"f800";
    tmp(27592) := x"f800";
    tmp(27593) := x"f800";
    tmp(27594) := x"f800";
    tmp(27595) := x"f800";
    tmp(27596) := x"f800";
    tmp(27597) := x"0840";
    tmp(27598) := x"0840";
    tmp(27599) := x"0840";
    tmp(27600) := x"0000";
    tmp(27601) := x"0022";
    tmp(27602) := x"0022";
    tmp(27603) := x"0022";
    tmp(27604) := x"0022";
    tmp(27605) := x"0022";
    tmp(27606) := x"0022";
    tmp(27607) := x"0021";
    tmp(27608) := x"0021";
    tmp(27609) := x"0022";
    tmp(27610) := x"0022";
    tmp(27611) := x"0022";
    tmp(27612) := x"0021";
    tmp(27613) := x"0842";
    tmp(27614) := x"0841";
    tmp(27615) := x"0821";
    tmp(27616) := x"0820";
    tmp(27617) := x"0021";
    tmp(27618) := x"0841";
    tmp(27619) := x"0041";
    tmp(27620) := x"0082";
    tmp(27621) := x"00a3";
    tmp(27622) := x"00a3";
    tmp(27623) := x"00a4";
    tmp(27624) := x"00a3";
    tmp(27625) := x"00a3";
    tmp(27626) := x"0083";
    tmp(27627) := x"00a4";
    tmp(27628) := x"00c4";
    tmp(27629) := x"08c4";
    tmp(27630) := x"08c4";
    tmp(27631) := x"08c4";
    tmp(27632) := x"08a4";
    tmp(27633) := x"08a3";
    tmp(27634) := x"08a3";
    tmp(27635) := x"08a4";
    tmp(27636) := x"08a3";
    tmp(27637) := x"08c4";
    tmp(27638) := x"08c3";
    tmp(27639) := x"08c4";
    tmp(27640) := x"08c4";
    tmp(27641) := x"08c4";
    tmp(27642) := x"08e4";
    tmp(27643) := x"08c4";
    tmp(27644) := x"08a3";
    tmp(27645) := x"08e4";
    tmp(27646) := x"08c4";
    tmp(27647) := x"0905";
    tmp(27648) := x"08e4";
    tmp(27649) := x"08a3";
    tmp(27650) := x"08c4";
    tmp(27651) := x"08e4";
    tmp(27652) := x"0904";
    tmp(27653) := x"0905";
    tmp(27654) := x"0905";
    tmp(27655) := x"0925";
    tmp(27656) := x"1167";
    tmp(27657) := x"1a29";
    tmp(27658) := x"0925";
    tmp(27659) := x"0925";
    tmp(27660) := x"0946";
    tmp(27661) := x"0967";
    tmp(27662) := x"0967";
    tmp(27663) := x"0967";
    tmp(27664) := x"0946";
    tmp(27665) := x"0967";
    tmp(27666) := x"0987";
    tmp(27667) := x"0946";
    tmp(27668) := x"0925";
    tmp(27669) := x"0925";
    tmp(27670) := x"0924";
    tmp(27671) := x"0924";
    tmp(27672) := x"0924";
    tmp(27673) := x"0945";
    tmp(27674) := x"0925";
    tmp(27675) := x"0905";
    tmp(27676) := x"0924";
    tmp(27677) := x"0925";
    tmp(27678) := x"0945";
    tmp(27679) := x"0965";
    tmp(27680) := x"1165";
    tmp(27681) := x"1186";
    tmp(27682) := x"1186";
    tmp(27683) := x"11a7";
    tmp(27684) := x"19e8";
    tmp(27685) := x"21e8";
    tmp(27686) := x"42ee";
    tmp(27687) := x"9537";
    tmp(27688) := x"df1f";
    tmp(27689) := x"f79f";
    tmp(27690) := x"ffff";
    tmp(27691) := x"ffff";
    tmp(27692) := x"ffff";
    tmp(27693) := x"ffff";
    tmp(27694) := x"ffff";
    tmp(27695) := x"ffff";
    tmp(27696) := x"ffff";
    tmp(27697) := x"ffff";
    tmp(27698) := x"ffff";
    tmp(27699) := x"ffff";
    tmp(27700) := x"ffff";
    tmp(27701) := x"ffff";
    tmp(27702) := x"ffff";
    tmp(27703) := x"ffff";
    tmp(27704) := x"ffff";
    tmp(27705) := x"ffff";
    tmp(27706) := x"ffff";
    tmp(27707) := x"ffff";
    tmp(27708) := x"ffff";
    tmp(27709) := x"f7fe";
    tmp(27710) := x"dfb9";
    tmp(27711) := x"be93";
    tmp(27712) := x"8d2d";
    tmp(27713) := x"6c09";
    tmp(27714) := x"4b05";
    tmp(27715) := x"2a22";
    tmp(27716) := x"1981";
    tmp(27717) := x"1140";
    tmp(27718) := x"1140";
    tmp(27719) := x"1981";
    tmp(27720) := x"1981";
    tmp(27721) := x"1961";
    tmp(27722) := x"1941";
    tmp(27723) := x"1121";
    tmp(27724) := x"1101";
    tmp(27725) := x"1101";
    tmp(27726) := x"1101";
    tmp(27727) := x"1121";
    tmp(27728) := x"2181";
    tmp(27729) := x"3a43";
    tmp(27730) := x"52e5";
    tmp(27731) := x"6b68";
    tmp(27732) := x"7bca";
    tmp(27733) := x"840c";
    tmp(27734) := x"8c8d";
    tmp(27735) := x"948e";
    tmp(27736) := x"946d";
    tmp(27737) := x"7baa";
    tmp(27738) := x"6b48";
    tmp(27739) := x"5ac6";
    tmp(27740) := x"4a44";
    tmp(27741) := x"39e3";
    tmp(27742) := x"2982";
    tmp(27743) := x"2141";
    tmp(27744) := x"1901";
    tmp(27745) := x"1901";
    tmp(27746) := x"1901";
    tmp(27747) := x"1921";
    tmp(27748) := x"2161";
    tmp(27749) := x"31a2";
    tmp(27750) := x"3a02";
    tmp(27751) := x"4a63";
    tmp(27752) := x"62e5";
    tmp(27753) := x"7367";
    tmp(27754) := x"93e9";
    tmp(27755) := x"acab";
    tmp(27756) := x"bd4c";
    tmp(27757) := x"bd4d";
    tmp(27758) := x"bd2d";
    tmp(27759) := x"bd2d";
    tmp(27760) := x"b4cc";
    tmp(27761) := x"ac8c";
    tmp(27762) := x"a46c";
    tmp(27763) := x"9c4b";
    tmp(27764) := x"940b";
    tmp(27765) := x"83ca";
    tmp(27766) := x"7369";
    tmp(27767) := x"7348";
    tmp(27768) := x"6b07";
    tmp(27769) := x"5ac7";
    tmp(27770) := x"5286";
    tmp(27771) := x"5266";
    tmp(27772) := x"5287";
    tmp(27773) := x"5aa7";
    tmp(27774) := x"5aa7";
    tmp(27775) := x"62c7";
    tmp(27776) := x"62c8";
    tmp(27777) := x"7329";
    tmp(27778) := x"836c";
    tmp(27779) := x"93ef";
    tmp(27780) := x"9c31";
    tmp(27781) := x"ac92";
    tmp(27782) := x"b4f4";
    tmp(27783) := x"b516";
    tmp(27784) := x"bd38";
    tmp(27785) := x"bd38";
    tmp(27786) := x"bd18";
    tmp(27787) := x"b4d8";
    tmp(27788) := x"b4b7";
    tmp(27789) := x"b4b7";
    tmp(27790) := x"b4b7";
    tmp(27791) := x"ac75";
    tmp(27792) := x"b4d6";
    tmp(27793) := x"b496";
    tmp(27794) := x"a434";
    tmp(27795) := x"a434";
    tmp(27796) := x"ac55";
    tmp(27797) := x"f800";
    tmp(27798) := x"f800";
    tmp(27799) := x"f800";
    tmp(27800) := x"f800";
    tmp(27801) := x"f800";
    tmp(27802) := x"f800";
    tmp(27803) := x"f800";
    tmp(27804) := x"f800";
    tmp(27805) := x"f800";
    tmp(27806) := x"f800";
    tmp(27807) := x"f800";
    tmp(27808) := x"f800";
    tmp(27809) := x"f800";
    tmp(27810) := x"f800";
    tmp(27811) := x"f800";
    tmp(27812) := x"f800";
    tmp(27813) := x"f800";
    tmp(27814) := x"f800";
    tmp(27815) := x"f800";
    tmp(27816) := x"f800";
    tmp(27817) := x"f800";
    tmp(27818) := x"f800";
    tmp(27819) := x"f800";
    tmp(27820) := x"f800";
    tmp(27821) := x"f800";
    tmp(27822) := x"f800";
    tmp(27823) := x"f800";
    tmp(27824) := x"f800";
    tmp(27825) := x"f800";
    tmp(27826) := x"f800";
    tmp(27827) := x"f800";
    tmp(27828) := x"f800";
    tmp(27829) := x"f800";
    tmp(27830) := x"f800";
    tmp(27831) := x"f800";
    tmp(27832) := x"f800";
    tmp(27833) := x"f800";
    tmp(27834) := x"f800";
    tmp(27835) := x"f800";
    tmp(27836) := x"f800";
    tmp(27837) := x"0840";
    tmp(27838) := x"0840";
    tmp(27839) := x"0840";
    tmp(27840) := x"0000";
    tmp(27841) := x"0000";
    tmp(27842) := x"0000";
    tmp(27843) := x"0020";
    tmp(27844) := x"0020";
    tmp(27845) := x"0020";
    tmp(27846) := x"0020";
    tmp(27847) := x"0020";
    tmp(27848) := x"0020";
    tmp(27849) := x"0020";
    tmp(27850) := x"0021";
    tmp(27851) := x"0021";
    tmp(27852) := x"0820";
    tmp(27853) := x"0821";
    tmp(27854) := x"0821";
    tmp(27855) := x"0821";
    tmp(27856) := x"0821";
    tmp(27857) := x"0020";
    tmp(27858) := x"0020";
    tmp(27859) := x"0020";
    tmp(27860) := x"0041";
    tmp(27861) := x"0062";
    tmp(27862) := x"00a3";
    tmp(27863) := x"00a3";
    tmp(27864) := x"00a3";
    tmp(27865) := x"0082";
    tmp(27866) := x"00a3";
    tmp(27867) := x"00c4";
    tmp(27868) := x"00c4";
    tmp(27869) := x"08c4";
    tmp(27870) := x"08e4";
    tmp(27871) := x"08c4";
    tmp(27872) := x"08c4";
    tmp(27873) := x"08c4";
    tmp(27874) := x"08c4";
    tmp(27875) := x"08a4";
    tmp(27876) := x"08c4";
    tmp(27877) := x"08e4";
    tmp(27878) := x"08e4";
    tmp(27879) := x"08e4";
    tmp(27880) := x"08e5";
    tmp(27881) := x"08c4";
    tmp(27882) := x"08a3";
    tmp(27883) := x"08a3";
    tmp(27884) := x"08a3";
    tmp(27885) := x"08e4";
    tmp(27886) := x"0904";
    tmp(27887) := x"0905";
    tmp(27888) := x"0925";
    tmp(27889) := x"0862";
    tmp(27890) := x"08c4";
    tmp(27891) := x"0905";
    tmp(27892) := x"0925";
    tmp(27893) := x"0925";
    tmp(27894) := x"1146";
    tmp(27895) := x"0925";
    tmp(27896) := x"0926";
    tmp(27897) := x"1187";
    tmp(27898) := x"1166";
    tmp(27899) := x"0966";
    tmp(27900) := x"0947";
    tmp(27901) := x"0967";
    tmp(27902) := x"0947";
    tmp(27903) := x"0947";
    tmp(27904) := x"0946";
    tmp(27905) := x"0926";
    tmp(27906) := x"0946";
    tmp(27907) := x"0946";
    tmp(27908) := x"0905";
    tmp(27909) := x"0905";
    tmp(27910) := x"0925";
    tmp(27911) := x"0925";
    tmp(27912) := x"0925";
    tmp(27913) := x"0966";
    tmp(27914) := x"0946";
    tmp(27915) := x"0946";
    tmp(27916) := x"0966";
    tmp(27917) := x"0966";
    tmp(27918) := x"11c8";
    tmp(27919) := x"1a29";
    tmp(27920) := x"19e8";
    tmp(27921) := x"1987";
    tmp(27922) := x"1987";
    tmp(27923) := x"3a8d";
    tmp(27924) := x"8cb6";
    tmp(27925) := x"df1e";
    tmp(27926) := x"ffff";
    tmp(27927) := x"ffff";
    tmp(27928) := x"ffff";
    tmp(27929) := x"ffff";
    tmp(27930) := x"ffff";
    tmp(27931) := x"ffff";
    tmp(27932) := x"ffff";
    tmp(27933) := x"ffff";
    tmp(27934) := x"ffff";
    tmp(27935) := x"ffff";
    tmp(27936) := x"ffff";
    tmp(27937) := x"ffff";
    tmp(27938) := x"ffff";
    tmp(27939) := x"ffff";
    tmp(27940) := x"ffff";
    tmp(27941) := x"ffff";
    tmp(27942) := x"ffff";
    tmp(27943) := x"ffff";
    tmp(27944) := x"ffff";
    tmp(27945) := x"ffff";
    tmp(27946) := x"ffff";
    tmp(27947) := x"f7ff";
    tmp(27948) := x"effe";
    tmp(27949) := x"d79a";
    tmp(27950) := x"be94";
    tmp(27951) := x"9d8f";
    tmp(27952) := x"746a";
    tmp(27953) := x"5346";
    tmp(27954) := x"3283";
    tmp(27955) := x"21c1";
    tmp(27956) := x"1140";
    tmp(27957) := x"1120";
    tmp(27958) := x"1140";
    tmp(27959) := x"1981";
    tmp(27960) := x"21a1";
    tmp(27961) := x"1981";
    tmp(27962) := x"1941";
    tmp(27963) := x"1121";
    tmp(27964) := x"1121";
    tmp(27965) := x"1121";
    tmp(27966) := x"1101";
    tmp(27967) := x"1101";
    tmp(27968) := x"1921";
    tmp(27969) := x"29a2";
    tmp(27970) := x"3a63";
    tmp(27971) := x"5306";
    tmp(27972) := x"6b88";
    tmp(27973) := x"73a9";
    tmp(27974) := x"7c0b";
    tmp(27975) := x"8c6c";
    tmp(27976) := x"8c4c";
    tmp(27977) := x"8c0c";
    tmp(27978) := x"7baa";
    tmp(27979) := x"6b07";
    tmp(27980) := x"5aa6";
    tmp(27981) := x"4a44";
    tmp(27982) := x"31c3";
    tmp(27983) := x"2982";
    tmp(27984) := x"2141";
    tmp(27985) := x"1921";
    tmp(27986) := x"1921";
    tmp(27987) := x"1921";
    tmp(27988) := x"2141";
    tmp(27989) := x"2161";
    tmp(27990) := x"29a2";
    tmp(27991) := x"3a02";
    tmp(27992) := x"4a63";
    tmp(27993) := x"62e5";
    tmp(27994) := x"7b47";
    tmp(27995) := x"9409";
    tmp(27996) := x"acab";
    tmp(27997) := x"accb";
    tmp(27998) := x"b50c";
    tmp(27999) := x"accb";
    tmp(28000) := x"accc";
    tmp(28001) := x"ac8c";
    tmp(28002) := x"b4cd";
    tmp(28003) := x"a46b";
    tmp(28004) := x"9c2b";
    tmp(28005) := x"8bca";
    tmp(28006) := x"83ca";
    tmp(28007) := x"7baa";
    tmp(28008) := x"6b48";
    tmp(28009) := x"62e7";
    tmp(28010) := x"5ac6";
    tmp(28011) := x"5286";
    tmp(28012) := x"5266";
    tmp(28013) := x"5267";
    tmp(28014) := x"5267";
    tmp(28015) := x"5266";
    tmp(28016) := x"62c8";
    tmp(28017) := x"6b09";
    tmp(28018) := x"7b4c";
    tmp(28019) := x"8bae";
    tmp(28020) := x"9c11";
    tmp(28021) := x"a493";
    tmp(28022) := x"acd4";
    tmp(28023) := x"acd5";
    tmp(28024) := x"b4f7";
    tmp(28025) := x"bcf8";
    tmp(28026) := x"b4f8";
    tmp(28027) := x"b4d7";
    tmp(28028) := x"b4b7";
    tmp(28029) := x"b4d7";
    tmp(28030) := x"ac96";
    tmp(28031) := x"ac75";
    tmp(28032) := x"ac95";
    tmp(28033) := x"ac55";
    tmp(28034) := x"a435";
    tmp(28035) := x"a415";
    tmp(28036) := x"a416";
    tmp(28037) := x"f800";
    tmp(28038) := x"f800";
    tmp(28039) := x"f800";
    tmp(28040) := x"f800";
    tmp(28041) := x"f800";
    tmp(28042) := x"f800";
    tmp(28043) := x"f800";
    tmp(28044) := x"f800";
    tmp(28045) := x"f800";
    tmp(28046) := x"f800";
    tmp(28047) := x"f800";
    tmp(28048) := x"f800";
    tmp(28049) := x"f800";
    tmp(28050) := x"f800";
    tmp(28051) := x"f800";
    tmp(28052) := x"f800";
    tmp(28053) := x"f800";
    tmp(28054) := x"f800";
    tmp(28055) := x"f800";
    tmp(28056) := x"f800";
    tmp(28057) := x"f800";
    tmp(28058) := x"f800";
    tmp(28059) := x"f800";
    tmp(28060) := x"f800";
    tmp(28061) := x"f800";
    tmp(28062) := x"f800";
    tmp(28063) := x"f800";
    tmp(28064) := x"f800";
    tmp(28065) := x"f800";
    tmp(28066) := x"f800";
    tmp(28067) := x"f800";
    tmp(28068) := x"f800";
    tmp(28069) := x"f800";
    tmp(28070) := x"f800";
    tmp(28071) := x"f800";
    tmp(28072) := x"f800";
    tmp(28073) := x"f800";
    tmp(28074) := x"f800";
    tmp(28075) := x"f800";
    tmp(28076) := x"f800";
    tmp(28077) := x"0840";
    tmp(28078) := x"0840";
    tmp(28079) := x"0840";
    tmp(28080) := x"0000";
    tmp(28081) := x"0000";
    tmp(28082) := x"0000";
    tmp(28083) := x"0000";
    tmp(28084) := x"0020";
    tmp(28085) := x"0020";
    tmp(28086) := x"0020";
    tmp(28087) := x"0020";
    tmp(28088) := x"0021";
    tmp(28089) := x"0020";
    tmp(28090) := x"0020";
    tmp(28091) := x"0020";
    tmp(28092) := x"0020";
    tmp(28093) := x"0020";
    tmp(28094) := x"0021";
    tmp(28095) := x"0020";
    tmp(28096) := x"0020";
    tmp(28097) := x"0021";
    tmp(28098) := x"0021";
    tmp(28099) := x"0020";
    tmp(28100) := x"0021";
    tmp(28101) := x"0041";
    tmp(28102) := x"0083";
    tmp(28103) := x"00a3";
    tmp(28104) := x"00a3";
    tmp(28105) := x"00a3";
    tmp(28106) := x"00a4";
    tmp(28107) := x"00c4";
    tmp(28108) := x"00c5";
    tmp(28109) := x"08c5";
    tmp(28110) := x"08e5";
    tmp(28111) := x"08e5";
    tmp(28112) := x"08e4";
    tmp(28113) := x"08c4";
    tmp(28114) := x"08a4";
    tmp(28115) := x"08c4";
    tmp(28116) := x"08c4";
    tmp(28117) := x"08c4";
    tmp(28118) := x"08c4";
    tmp(28119) := x"08c4";
    tmp(28120) := x"08c4";
    tmp(28121) := x"08c4";
    tmp(28122) := x"08c3";
    tmp(28123) := x"08c4";
    tmp(28124) := x"08e4";
    tmp(28125) := x"08e5";
    tmp(28126) := x"08e4";
    tmp(28127) := x"08e4";
    tmp(28128) := x"0905";
    tmp(28129) := x"08a3";
    tmp(28130) := x"0926";
    tmp(28131) := x"0925";
    tmp(28132) := x"08e4";
    tmp(28133) := x"0905";
    tmp(28134) := x"1146";
    tmp(28135) := x"1146";
    tmp(28136) := x"0905";
    tmp(28137) := x"08a3";
    tmp(28138) := x"19c8";
    tmp(28139) := x"08c3";
    tmp(28140) := x"0966";
    tmp(28141) := x"0926";
    tmp(28142) := x"0927";
    tmp(28143) := x"0927";
    tmp(28144) := x"0926";
    tmp(28145) := x"0925";
    tmp(28146) := x"0946";
    tmp(28147) := x"0946";
    tmp(28148) := x"0905";
    tmp(28149) := x"0905";
    tmp(28150) := x"0946";
    tmp(28151) := x"0966";
    tmp(28152) := x"0966";
    tmp(28153) := x"0966";
    tmp(28154) := x"09a8";
    tmp(28155) := x"11e9";
    tmp(28156) := x"124a";
    tmp(28157) := x"1229";
    tmp(28158) := x"1a2a";
    tmp(28159) := x"224b";
    tmp(28160) := x"4b2f";
    tmp(28161) := x"9d38";
    tmp(28162) := x"f79f";
    tmp(28163) := x"ffff";
    tmp(28164) := x"ffff";
    tmp(28165) := x"ffff";
    tmp(28166) := x"ffff";
    tmp(28167) := x"ffff";
    tmp(28168) := x"ffff";
    tmp(28169) := x"ffff";
    tmp(28170) := x"ffff";
    tmp(28171) := x"ffff";
    tmp(28172) := x"ffff";
    tmp(28173) := x"ffff";
    tmp(28174) := x"ffff";
    tmp(28175) := x"ffff";
    tmp(28176) := x"ffff";
    tmp(28177) := x"ffff";
    tmp(28178) := x"ffff";
    tmp(28179) := x"ffff";
    tmp(28180) := x"ffff";
    tmp(28181) := x"ffff";
    tmp(28182) := x"ffff";
    tmp(28183) := x"ffff";
    tmp(28184) := x"ffff";
    tmp(28185) := x"f7ff";
    tmp(28186) := x"efdf";
    tmp(28187) := x"d79d";
    tmp(28188) := x"cf19";
    tmp(28189) := x"beb6";
    tmp(28190) := x"a5d1";
    tmp(28191) := x"7c6b";
    tmp(28192) := x"5b87";
    tmp(28193) := x"3ac4";
    tmp(28194) := x"2a02";
    tmp(28195) := x"1161";
    tmp(28196) := x"0920";
    tmp(28197) := x"0920";
    tmp(28198) := x"1161";
    tmp(28199) := x"19a1";
    tmp(28200) := x"21c1";
    tmp(28201) := x"21a1";
    tmp(28202) := x"1961";
    tmp(28203) := x"1941";
    tmp(28204) := x"1921";
    tmp(28205) := x"1121";
    tmp(28206) := x"1101";
    tmp(28207) := x"1101";
    tmp(28208) := x"1101";
    tmp(28209) := x"1961";
    tmp(28210) := x"29e2";
    tmp(28211) := x"4264";
    tmp(28212) := x"5b06";
    tmp(28213) := x"6b88";
    tmp(28214) := x"73c9";
    tmp(28215) := x"7c0a";
    tmp(28216) := x"844b";
    tmp(28217) := x"840b";
    tmp(28218) := x"83ea";
    tmp(28219) := x"7369";
    tmp(28220) := x"62e7";
    tmp(28221) := x"5285";
    tmp(28222) := x"4224";
    tmp(28223) := x"31c3";
    tmp(28224) := x"2982";
    tmp(28225) := x"2141";
    tmp(28226) := x"1921";
    tmp(28227) := x"1921";
    tmp(28228) := x"2141";
    tmp(28229) := x"2141";
    tmp(28230) := x"2161";
    tmp(28231) := x"31a2";
    tmp(28232) := x"4202";
    tmp(28233) := x"5263";
    tmp(28234) := x"62c5";
    tmp(28235) := x"7b67";
    tmp(28236) := x"93e9";
    tmp(28237) := x"a48b";
    tmp(28238) := x"b4ec";
    tmp(28239) := x"accc";
    tmp(28240) := x"a48c";
    tmp(28241) := x"a48b";
    tmp(28242) := x"a46b";
    tmp(28243) := x"940b";
    tmp(28244) := x"9c0b";
    tmp(28245) := x"940b";
    tmp(28246) := x"8baa";
    tmp(28247) := x"7349";
    tmp(28248) := x"6b48";
    tmp(28249) := x"6ae7";
    tmp(28250) := x"5ac7";
    tmp(28251) := x"5286";
    tmp(28252) := x"5246";
    tmp(28253) := x"4a46";
    tmp(28254) := x"5246";
    tmp(28255) := x"5246";
    tmp(28256) := x"5a87";
    tmp(28257) := x"6b09";
    tmp(28258) := x"7b4b";
    tmp(28259) := x"93ce";
    tmp(28260) := x"93f0";
    tmp(28261) := x"a472";
    tmp(28262) := x"ac95";
    tmp(28263) := x"b4d5";
    tmp(28264) := x"b4d6";
    tmp(28265) := x"b4d7";
    tmp(28266) := x"acb7";
    tmp(28267) := x"acb7";
    tmp(28268) := x"ac97";
    tmp(28269) := x"a495";
    tmp(28270) := x"ac76";
    tmp(28271) := x"ac76";
    tmp(28272) := x"ac95";
    tmp(28273) := x"ac55";
    tmp(28274) := x"a454";
    tmp(28275) := x"9c14";
    tmp(28276) := x"a415";
    tmp(28277) := x"f800";
    tmp(28278) := x"f800";
    tmp(28279) := x"f800";
    tmp(28280) := x"f800";
    tmp(28281) := x"f800";
    tmp(28282) := x"f800";
    tmp(28283) := x"f800";
    tmp(28284) := x"f800";
    tmp(28285) := x"f800";
    tmp(28286) := x"f800";
    tmp(28287) := x"f800";
    tmp(28288) := x"f800";
    tmp(28289) := x"f800";
    tmp(28290) := x"f800";
    tmp(28291) := x"f800";
    tmp(28292) := x"f800";
    tmp(28293) := x"f800";
    tmp(28294) := x"f800";
    tmp(28295) := x"f800";
    tmp(28296) := x"f800";
    tmp(28297) := x"f800";
    tmp(28298) := x"f800";
    tmp(28299) := x"f800";
    tmp(28300) := x"f800";
    tmp(28301) := x"f800";
    tmp(28302) := x"f800";
    tmp(28303) := x"f800";
    tmp(28304) := x"f800";
    tmp(28305) := x"f800";
    tmp(28306) := x"f800";
    tmp(28307) := x"f800";
    tmp(28308) := x"f800";
    tmp(28309) := x"f800";
    tmp(28310) := x"f800";
    tmp(28311) := x"f800";
    tmp(28312) := x"f800";
    tmp(28313) := x"f800";
    tmp(28314) := x"f800";
    tmp(28315) := x"f800";
    tmp(28316) := x"f800";
    tmp(28317) := x"0840";
    tmp(28318) := x"0840";
    tmp(28319) := x"0840";
    tmp(28320) := x"0000";
    tmp(28321) := x"0021";
    tmp(28322) := x"0021";
    tmp(28323) := x"0000";
    tmp(28324) := x"0000";
    tmp(28325) := x"0020";
    tmp(28326) := x"0021";
    tmp(28327) := x"0021";
    tmp(28328) := x"0021";
    tmp(28329) := x"0021";
    tmp(28330) := x"0021";
    tmp(28331) := x"0021";
    tmp(28332) := x"0021";
    tmp(28333) := x"0020";
    tmp(28334) := x"0020";
    tmp(28335) := x"0021";
    tmp(28336) := x"0021";
    tmp(28337) := x"0021";
    tmp(28338) := x"0841";
    tmp(28339) := x"0021";
    tmp(28340) := x"0041";
    tmp(28341) := x"0062";
    tmp(28342) := x"0083";
    tmp(28343) := x"00a4";
    tmp(28344) := x"08c4";
    tmp(28345) := x"00c4";
    tmp(28346) := x"08e5";
    tmp(28347) := x"08e5";
    tmp(28348) := x"0906";
    tmp(28349) := x"0906";
    tmp(28350) := x"0905";
    tmp(28351) := x"08e5";
    tmp(28352) := x"0905";
    tmp(28353) := x"08e5";
    tmp(28354) := x"08c4";
    tmp(28355) := x"08c4";
    tmp(28356) := x"08e4";
    tmp(28357) := x"08e4";
    tmp(28358) := x"08e5";
    tmp(28359) := x"08e5";
    tmp(28360) := x"08e4";
    tmp(28361) := x"08c4";
    tmp(28362) := x"08c4";
    tmp(28363) := x"08e4";
    tmp(28364) := x"08e4";
    tmp(28365) := x"08e4";
    tmp(28366) := x"08e4";
    tmp(28367) := x"08e4";
    tmp(28368) := x"08c3";
    tmp(28369) := x"08c4";
    tmp(28370) := x"0905";
    tmp(28371) := x"08e4";
    tmp(28372) := x"0904";
    tmp(28373) := x"08e4";
    tmp(28374) := x"10e3";
    tmp(28375) := x"08c3";
    tmp(28376) := x"0904";
    tmp(28377) := x"08c3";
    tmp(28378) := x"1187";
    tmp(28379) := x"1165";
    tmp(28380) := x"08e2";
    tmp(28381) := x"1187";
    tmp(28382) := x"0968";
    tmp(28383) := x"0926";
    tmp(28384) := x"0926";
    tmp(28385) := x"0946";
    tmp(28386) := x"0925";
    tmp(28387) := x"0905";
    tmp(28388) := x"0925";
    tmp(28389) := x"0946";
    tmp(28390) := x"0966";
    tmp(28391) := x"0967";
    tmp(28392) := x"09a7";
    tmp(28393) := x"122a";
    tmp(28394) := x"126c";
    tmp(28395) := x"1aac";
    tmp(28396) := x"1a6b";
    tmp(28397) := x"2a8c";
    tmp(28398) := x"5bb1";
    tmp(28399) := x"add9";
    tmp(28400) := x"ffff";
    tmp(28401) := x"ffff";
    tmp(28402) := x"ffff";
    tmp(28403) := x"ffff";
    tmp(28404) := x"ffff";
    tmp(28405) := x"ffff";
    tmp(28406) := x"ffff";
    tmp(28407) := x"ffff";
    tmp(28408) := x"ffff";
    tmp(28409) := x"ffff";
    tmp(28410) := x"ffff";
    tmp(28411) := x"ffff";
    tmp(28412) := x"ffff";
    tmp(28413) := x"ffff";
    tmp(28414) := x"ffff";
    tmp(28415) := x"ffff";
    tmp(28416) := x"ffff";
    tmp(28417) := x"ffff";
    tmp(28418) := x"ffff";
    tmp(28419) := x"ffff";
    tmp(28420) := x"ffff";
    tmp(28421) := x"ffff";
    tmp(28422) := x"ffff";
    tmp(28423) := x"efff";
    tmp(28424) := x"efdf";
    tmp(28425) := x"d79f";
    tmp(28426) := x"c71c";
    tmp(28427) := x"cf1a";
    tmp(28428) := x"b654";
    tmp(28429) := x"9db1";
    tmp(28430) := x"7c8c";
    tmp(28431) := x"5ba8";
    tmp(28432) := x"42e5";
    tmp(28433) := x"3243";
    tmp(28434) := x"19a1";
    tmp(28435) := x"1141";
    tmp(28436) := x"0900";
    tmp(28437) := x"1120";
    tmp(28438) := x"1961";
    tmp(28439) := x"19a1";
    tmp(28440) := x"21c1";
    tmp(28441) := x"21c1";
    tmp(28442) := x"1981";
    tmp(28443) := x"1941";
    tmp(28444) := x"1921";
    tmp(28445) := x"1121";
    tmp(28446) := x"1101";
    tmp(28447) := x"1101";
    tmp(28448) := x"1121";
    tmp(28449) := x"1121";
    tmp(28450) := x"2161";
    tmp(28451) := x"31e2";
    tmp(28452) := x"4284";
    tmp(28453) := x"5306";
    tmp(28454) := x"6b87";
    tmp(28455) := x"73a9";
    tmp(28456) := x"73ca";
    tmp(28457) := x"83ea";
    tmp(28458) := x"83ca";
    tmp(28459) := x"7bc9";
    tmp(28460) := x"6b48";
    tmp(28461) := x"62e6";
    tmp(28462) := x"5285";
    tmp(28463) := x"4224";
    tmp(28464) := x"31c3";
    tmp(28465) := x"2962";
    tmp(28466) := x"2121";
    tmp(28467) := x"1921";
    tmp(28468) := x"1921";
    tmp(28469) := x"2141";
    tmp(28470) := x"2141";
    tmp(28471) := x"2161";
    tmp(28472) := x"2981";
    tmp(28473) := x"39e2";
    tmp(28474) := x"4a64";
    tmp(28475) := x"62e5";
    tmp(28476) := x"7b67";
    tmp(28477) := x"942a";
    tmp(28478) := x"a48b";
    tmp(28479) := x"a46b";
    tmp(28480) := x"9c4b";
    tmp(28481) := x"942a";
    tmp(28482) := x"940b";
    tmp(28483) := x"93ea";
    tmp(28484) := x"8bca";
    tmp(28485) := x"8bca";
    tmp(28486) := x"83aa";
    tmp(28487) := x"7b69";
    tmp(28488) := x"7348";
    tmp(28489) := x"6307";
    tmp(28490) := x"5aa7";
    tmp(28491) := x"5266";
    tmp(28492) := x"5246";
    tmp(28493) := x"4a25";
    tmp(28494) := x"4a25";
    tmp(28495) := x"5246";
    tmp(28496) := x"5a87";
    tmp(28497) := x"6b0a";
    tmp(28498) := x"7b6c";
    tmp(28499) := x"8bad";
    tmp(28500) := x"9410";
    tmp(28501) := x"9c12";
    tmp(28502) := x"a453";
    tmp(28503) := x"a474";
    tmp(28504) := x"acb6";
    tmp(28505) := x"b4d7";
    tmp(28506) := x"b4d7";
    tmp(28507) := x"b4d7";
    tmp(28508) := x"b4d7";
    tmp(28509) := x"a476";
    tmp(28510) := x"ac77";
    tmp(28511) := x"ac76";
    tmp(28512) := x"ac75";
    tmp(28513) := x"ac75";
    tmp(28514) := x"a434";
    tmp(28515) := x"9c15";
    tmp(28516) := x"9c15";
    tmp(28517) := x"f800";
    tmp(28518) := x"f800";
    tmp(28519) := x"f800";
    tmp(28520) := x"f800";
    tmp(28521) := x"f800";
    tmp(28522) := x"f800";
    tmp(28523) := x"f800";
    tmp(28524) := x"f800";
    tmp(28525) := x"f800";
    tmp(28526) := x"f800";
    tmp(28527) := x"f800";
    tmp(28528) := x"f800";
    tmp(28529) := x"f800";
    tmp(28530) := x"f800";
    tmp(28531) := x"f800";
    tmp(28532) := x"f800";
    tmp(28533) := x"f800";
    tmp(28534) := x"f800";
    tmp(28535) := x"f800";
    tmp(28536) := x"f800";
    tmp(28537) := x"f800";
    tmp(28538) := x"f800";
    tmp(28539) := x"f800";
    tmp(28540) := x"f800";
    tmp(28541) := x"f800";
    tmp(28542) := x"f800";
    tmp(28543) := x"f800";
    tmp(28544) := x"f800";
    tmp(28545) := x"f800";
    tmp(28546) := x"f800";
    tmp(28547) := x"f800";
    tmp(28548) := x"f800";
    tmp(28549) := x"f800";
    tmp(28550) := x"f800";
    tmp(28551) := x"f800";
    tmp(28552) := x"f800";
    tmp(28553) := x"f800";
    tmp(28554) := x"f800";
    tmp(28555) := x"f800";
    tmp(28556) := x"f800";
    tmp(28557) := x"0840";
    tmp(28558) := x"0840";
    tmp(28559) := x"0840";
    tmp(28560) := x"0000";
    tmp(28561) := x"0021";
    tmp(28562) := x"0041";
    tmp(28563) := x"0021";
    tmp(28564) := x"0021";
    tmp(28565) := x"0041";
    tmp(28566) := x"0021";
    tmp(28567) := x"0021";
    tmp(28568) := x"0021";
    tmp(28569) := x"0020";
    tmp(28570) := x"0021";
    tmp(28571) := x"0041";
    tmp(28572) := x"0021";
    tmp(28573) := x"0021";
    tmp(28574) := x"0021";
    tmp(28575) := x"0041";
    tmp(28576) := x"0041";
    tmp(28577) := x"0021";
    tmp(28578) := x"0041";
    tmp(28579) := x"0021";
    tmp(28580) := x"0041";
    tmp(28581) := x"0042";
    tmp(28582) := x"0062";
    tmp(28583) := x"0083";
    tmp(28584) := x"00a3";
    tmp(28585) := x"00a3";
    tmp(28586) := x"00c4";
    tmp(28587) := x"08e5";
    tmp(28588) := x"08e5";
    tmp(28589) := x"08e5";
    tmp(28590) := x"08e5";
    tmp(28591) := x"08e5";
    tmp(28592) := x"08c4";
    tmp(28593) := x"08c4";
    tmp(28594) := x"00a4";
    tmp(28595) := x"08c4";
    tmp(28596) := x"08c4";
    tmp(28597) := x"0905";
    tmp(28598) := x"08e5";
    tmp(28599) := x"08a4";
    tmp(28600) := x"08c4";
    tmp(28601) := x"08c4";
    tmp(28602) := x"08c4";
    tmp(28603) := x"08e4";
    tmp(28604) := x"08e4";
    tmp(28605) := x"08e5";
    tmp(28606) := x"08c4";
    tmp(28607) := x"08e4";
    tmp(28608) := x"08e4";
    tmp(28609) := x"08e4";
    tmp(28610) := x"08e4";
    tmp(28611) := x"08e4";
    tmp(28612) := x"08e4";
    tmp(28613) := x"08a2";
    tmp(28614) := x"0841";
    tmp(28615) := x"0861";
    tmp(28616) := x"1105";
    tmp(28617) := x"08c4";
    tmp(28618) := x"0905";
    tmp(28619) := x"19e8";
    tmp(28620) := x"0861";
    tmp(28621) := x"1165";
    tmp(28622) := x"0905";
    tmp(28623) := x"08a3";
    tmp(28624) := x"0904";
    tmp(28625) := x"0966";
    tmp(28626) := x"0946";
    tmp(28627) := x"0925";
    tmp(28628) := x"0966";
    tmp(28629) := x"0987";
    tmp(28630) := x"0987";
    tmp(28631) := x"0987";
    tmp(28632) := x"120a";
    tmp(28633) := x"126b";
    tmp(28634) := x"1a6b";
    tmp(28635) := x"2a8b";
    tmp(28636) := x"534f";
    tmp(28637) := x"add7";
    tmp(28638) := x"ef1d";
    tmp(28639) := x"ff5d";
    tmp(28640) := x"ef1e";
    tmp(28641) := x"ff9f";
    tmp(28642) := x"ffbf";
    tmp(28643) := x"ffdf";
    tmp(28644) := x"ffdf";
    tmp(28645) := x"ffdf";
    tmp(28646) := x"ffff";
    tmp(28647) := x"ffff";
    tmp(28648) := x"ffff";
    tmp(28649) := x"ffff";
    tmp(28650) := x"ffff";
    tmp(28651) := x"ffff";
    tmp(28652) := x"ffff";
    tmp(28653) := x"ffff";
    tmp(28654) := x"ffff";
    tmp(28655) := x"ffff";
    tmp(28656) := x"ffff";
    tmp(28657) := x"ffff";
    tmp(28658) := x"ffff";
    tmp(28659) := x"ffff";
    tmp(28660) := x"ffff";
    tmp(28661) := x"f7df";
    tmp(28662) := x"efdf";
    tmp(28663) := x"d79f";
    tmp(28664) := x"cf3f";
    tmp(28665) := x"bedd";
    tmp(28666) := x"be99";
    tmp(28667) := x"ae36";
    tmp(28668) := x"9d72";
    tmp(28669) := x"84ad";
    tmp(28670) := x"6be9";
    tmp(28671) := x"4b26";
    tmp(28672) := x"3264";
    tmp(28673) := x"21c2";
    tmp(28674) := x"1161";
    tmp(28675) := x"1121";
    tmp(28676) := x"0900";
    tmp(28677) := x"1121";
    tmp(28678) := x"1981";
    tmp(28679) := x"21a1";
    tmp(28680) := x"21a1";
    tmp(28681) := x"21a1";
    tmp(28682) := x"1981";
    tmp(28683) := x"1961";
    tmp(28684) := x"1941";
    tmp(28685) := x"1121";
    tmp(28686) := x"1921";
    tmp(28687) := x"1121";
    tmp(28688) := x"1121";
    tmp(28689) := x"1101";
    tmp(28690) := x"1921";
    tmp(28691) := x"2181";
    tmp(28692) := x"3222";
    tmp(28693) := x"4a84";
    tmp(28694) := x"5b46";
    tmp(28695) := x"6b67";
    tmp(28696) := x"7388";
    tmp(28697) := x"7bc9";
    tmp(28698) := x"7be9";
    tmp(28699) := x"7ba8";
    tmp(28700) := x"7b89";
    tmp(28701) := x"7348";
    tmp(28702) := x"5ac6";
    tmp(28703) := x"5265";
    tmp(28704) := x"4224";
    tmp(28705) := x"31c3";
    tmp(28706) := x"2162";
    tmp(28707) := x"1921";
    tmp(28708) := x"1921";
    tmp(28709) := x"2121";
    tmp(28710) := x"2141";
    tmp(28711) := x"2161";
    tmp(28712) := x"2141";
    tmp(28713) := x"29a2";
    tmp(28714) := x"3a02";
    tmp(28715) := x"4a64";
    tmp(28716) := x"62e5";
    tmp(28717) := x"7b67";
    tmp(28718) := x"93e9";
    tmp(28719) := x"9c4a";
    tmp(28720) := x"9c4b";
    tmp(28721) := x"940a";
    tmp(28722) := x"93ea";
    tmp(28723) := x"8baa";
    tmp(28724) := x"8389";
    tmp(28725) := x"7b68";
    tmp(28726) := x"7b69";
    tmp(28727) := x"7b49";
    tmp(28728) := x"6b08";
    tmp(28729) := x"62c7";
    tmp(28730) := x"5aa7";
    tmp(28731) := x"5286";
    tmp(28732) := x"4a45";
    tmp(28733) := x"4205";
    tmp(28734) := x"4a05";
    tmp(28735) := x"5246";
    tmp(28736) := x"5a88";
    tmp(28737) := x"6aea";
    tmp(28738) := x"732b";
    tmp(28739) := x"8b8d";
    tmp(28740) := x"836e";
    tmp(28741) := x"93d1";
    tmp(28742) := x"9c11";
    tmp(28743) := x"93f2";
    tmp(28744) := x"a434";
    tmp(28745) := x"ac55";
    tmp(28746) := x"ac96";
    tmp(28747) := x"acb6";
    tmp(28748) := x"ac96";
    tmp(28749) := x"ac96";
    tmp(28750) := x"ac76";
    tmp(28751) := x"ac76";
    tmp(28752) := x"a455";
    tmp(28753) := x"a414";
    tmp(28754) := x"a456";
    tmp(28755) := x"9c15";
    tmp(28756) := x"9bf5";
    tmp(28757) := x"f800";
    tmp(28758) := x"f800";
    tmp(28759) := x"f800";
    tmp(28760) := x"f800";
    tmp(28761) := x"f800";
    tmp(28762) := x"f800";
    tmp(28763) := x"f800";
    tmp(28764) := x"f800";
    tmp(28765) := x"f800";
    tmp(28766) := x"f800";
    tmp(28767) := x"f800";
    tmp(28768) := x"f800";
    tmp(28769) := x"f800";
    tmp(28770) := x"f800";
    tmp(28771) := x"f800";
    tmp(28772) := x"f800";
    tmp(28773) := x"f800";
    tmp(28774) := x"f800";
    tmp(28775) := x"f800";
    tmp(28776) := x"f800";
    tmp(28777) := x"f800";
    tmp(28778) := x"f800";
    tmp(28779) := x"f800";
    tmp(28780) := x"f800";
    tmp(28781) := x"f800";
    tmp(28782) := x"f800";
    tmp(28783) := x"f800";
    tmp(28784) := x"f800";
    tmp(28785) := x"f800";
    tmp(28786) := x"f800";
    tmp(28787) := x"f800";
    tmp(28788) := x"f800";
    tmp(28789) := x"f800";
    tmp(28790) := x"f800";
    tmp(28791) := x"f800";
    tmp(28792) := x"f800";
    tmp(28793) := x"f800";
    tmp(28794) := x"f800";
    tmp(28795) := x"f800";
    tmp(28796) := x"f800";
    tmp(28797) := x"0840";
    tmp(28798) := x"0840";
    tmp(28799) := x"0840";
    tmp(28800) := x"0000";
    tmp(28801) := x"0021";
    tmp(28802) := x"0041";
    tmp(28803) := x"0021";
    tmp(28804) := x"0041";
    tmp(28805) := x"0041";
    tmp(28806) := x"0041";
    tmp(28807) := x"0041";
    tmp(28808) := x"0041";
    tmp(28809) := x"0042";
    tmp(28810) := x"0082";
    tmp(28811) := x"0083";
    tmp(28812) := x"0083";
    tmp(28813) := x"0083";
    tmp(28814) := x"0082";
    tmp(28815) := x"08a3";
    tmp(28816) := x"08a3";
    tmp(28817) := x"0882";
    tmp(28818) := x"0842";
    tmp(28819) := x"0021";
    tmp(28820) := x"0021";
    tmp(28821) := x"0020";
    tmp(28822) := x"0021";
    tmp(28823) := x"0062";
    tmp(28824) := x"00a3";
    tmp(28825) := x"00a3";
    tmp(28826) := x"00a3";
    tmp(28827) := x"00a4";
    tmp(28828) := x"00c4";
    tmp(28829) := x"08c4";
    tmp(28830) := x"08c4";
    tmp(28831) := x"08c4";
    tmp(28832) := x"08c4";
    tmp(28833) := x"08a4";
    tmp(28834) := x"00a4";
    tmp(28835) := x"08c4";
    tmp(28836) := x"08e5";
    tmp(28837) := x"08e4";
    tmp(28838) := x"08c4";
    tmp(28839) := x"08a3";
    tmp(28840) := x"08c3";
    tmp(28841) := x"08a3";
    tmp(28842) := x"08c4";
    tmp(28843) := x"08c4";
    tmp(28844) := x"08c4";
    tmp(28845) := x"08c4";
    tmp(28846) := x"08c4";
    tmp(28847) := x"08c4";
    tmp(28848) := x"08a3";
    tmp(28849) := x"08e4";
    tmp(28850) := x"0904";
    tmp(28851) := x"0904";
    tmp(28852) := x"0903";
    tmp(28853) := x"0882";
    tmp(28854) := x"0861";
    tmp(28855) := x"08c3";
    tmp(28856) := x"1125";
    tmp(28857) := x"1146";
    tmp(28858) := x"0904";
    tmp(28859) := x"1125";
    tmp(28860) := x"08a2";
    tmp(28861) := x"0861";
    tmp(28862) := x"0881";
    tmp(28863) := x"08a2";
    tmp(28864) := x"0925";
    tmp(28865) := x"0946";
    tmp(28866) := x"0966";
    tmp(28867) := x"09a8";
    tmp(28868) := x"0a0a";
    tmp(28869) := x"124b";
    tmp(28870) := x"122a";
    tmp(28871) := x"1209";
    tmp(28872) := x"1a29";
    tmp(28873) := x"2a49";
    tmp(28874) := x"4aeb";
    tmp(28875) := x"9491";
    tmp(28876) := x"c5b5";
    tmp(28877) := x"cdf6";
    tmp(28878) := x"ce18";
    tmp(28879) := x"e67b";
    tmp(28880) := x"eebc";
    tmp(28881) := x"eefe";
    tmp(28882) := x"f73f";
    tmp(28883) := x"f77f";
    tmp(28884) := x"ff9f";
    tmp(28885) := x"ffbf";
    tmp(28886) := x"ffbf";
    tmp(28887) := x"ffdf";
    tmp(28888) := x"ffff";
    tmp(28889) := x"ffff";
    tmp(28890) := x"ffff";
    tmp(28891) := x"ffff";
    tmp(28892) := x"ffff";
    tmp(28893) := x"ffdf";
    tmp(28894) := x"f7ff";
    tmp(28895) := x"efdf";
    tmp(28896) := x"f7df";
    tmp(28897) := x"efdf";
    tmp(28898) := x"efdf";
    tmp(28899) := x"e7bf";
    tmp(28900) := x"dfbf";
    tmp(28901) := x"d79f";
    tmp(28902) := x"cf5f";
    tmp(28903) := x"bede";
    tmp(28904) := x"b67c";
    tmp(28905) := x"a5f8";
    tmp(28906) := x"adf5";
    tmp(28907) := x"9d32";
    tmp(28908) := x"848e";
    tmp(28909) := x"6bea";
    tmp(28910) := x"5347";
    tmp(28911) := x"3aa5";
    tmp(28912) := x"2a03";
    tmp(28913) := x"1981";
    tmp(28914) := x"1141";
    tmp(28915) := x"1121";
    tmp(28916) := x"1121";
    tmp(28917) := x"1141";
    tmp(28918) := x"1981";
    tmp(28919) := x"21c1";
    tmp(28920) := x"21c1";
    tmp(28921) := x"1961";
    tmp(28922) := x"1961";
    tmp(28923) := x"1961";
    tmp(28924) := x"1941";
    tmp(28925) := x"1921";
    tmp(28926) := x"1921";
    tmp(28927) := x"1921";
    tmp(28928) := x"1921";
    tmp(28929) := x"1121";
    tmp(28930) := x"1121";
    tmp(28931) := x"1941";
    tmp(28932) := x"21a1";
    tmp(28933) := x"3a22";
    tmp(28934) := x"4aa4";
    tmp(28935) := x"6326";
    tmp(28936) := x"6b47";
    tmp(28937) := x"6b68";
    tmp(28938) := x"7388";
    tmp(28939) := x"7388";
    tmp(28940) := x"7b88";
    tmp(28941) := x"7368";
    tmp(28942) := x"6b27";
    tmp(28943) := x"5ac6";
    tmp(28944) := x"4a45";
    tmp(28945) := x"39e3";
    tmp(28946) := x"31a3";
    tmp(28947) := x"2162";
    tmp(28948) := x"2121";
    tmp(28949) := x"1921";
    tmp(28950) := x"2121";
    tmp(28951) := x"2141";
    tmp(28952) := x"2141";
    tmp(28953) := x"2161";
    tmp(28954) := x"31a2";
    tmp(28955) := x"39e2";
    tmp(28956) := x"4a64";
    tmp(28957) := x"62c5";
    tmp(28958) := x"7b67";
    tmp(28959) := x"8be9";
    tmp(28960) := x"940a";
    tmp(28961) := x"8bea";
    tmp(28962) := x"8bea";
    tmp(28963) := x"8389";
    tmp(28964) := x"8389";
    tmp(28965) := x"7347";
    tmp(28966) := x"7327";
    tmp(28967) := x"6b07";
    tmp(28968) := x"62c7";
    tmp(28969) := x"5aa6";
    tmp(28970) := x"5286";
    tmp(28971) := x"5266";
    tmp(28972) := x"4a45";
    tmp(28973) := x"4205";
    tmp(28974) := x"4a05";
    tmp(28975) := x"5246";
    tmp(28976) := x"5a87";
    tmp(28977) := x"62ca";
    tmp(28978) := x"6aea";
    tmp(28979) := x"7b4c";
    tmp(28980) := x"836d";
    tmp(28981) := x"836f";
    tmp(28982) := x"8bb0";
    tmp(28983) := x"8bb1";
    tmp(28984) := x"93d2";
    tmp(28985) := x"a415";
    tmp(28986) := x"ac76";
    tmp(28987) := x"ac96";
    tmp(28988) := x"ac97";
    tmp(28989) := x"ac96";
    tmp(28990) := x"ac76";
    tmp(28991) := x"ac76";
    tmp(28992) := x"a456";
    tmp(28993) := x"a415";
    tmp(28994) := x"a415";
    tmp(28995) := x"a456";
    tmp(28996) := x"9c15";
    tmp(28997) := x"f800";
    tmp(28998) := x"f800";
    tmp(28999) := x"f800";
    tmp(29000) := x"f800";
    tmp(29001) := x"f800";
    tmp(29002) := x"f800";
    tmp(29003) := x"f800";
    tmp(29004) := x"f800";
    tmp(29005) := x"f800";
    tmp(29006) := x"f800";
    tmp(29007) := x"f800";
    tmp(29008) := x"f800";
    tmp(29009) := x"f800";
    tmp(29010) := x"f800";
    tmp(29011) := x"f800";
    tmp(29012) := x"f800";
    tmp(29013) := x"f800";
    tmp(29014) := x"f800";
    tmp(29015) := x"f800";
    tmp(29016) := x"f800";
    tmp(29017) := x"f800";
    tmp(29018) := x"f800";
    tmp(29019) := x"f800";
    tmp(29020) := x"f800";
    tmp(29021) := x"f800";
    tmp(29022) := x"f800";
    tmp(29023) := x"f800";
    tmp(29024) := x"f800";
    tmp(29025) := x"f800";
    tmp(29026) := x"f800";
    tmp(29027) := x"f800";
    tmp(29028) := x"f800";
    tmp(29029) := x"f800";
    tmp(29030) := x"f800";
    tmp(29031) := x"f800";
    tmp(29032) := x"f800";
    tmp(29033) := x"f800";
    tmp(29034) := x"f800";
    tmp(29035) := x"f800";
    tmp(29036) := x"f800";
    tmp(29037) := x"0840";
    tmp(29038) := x"0840";
    tmp(29039) := x"0840";
    tmp(29040) := x"0000";
    tmp(29041) := x"0062";
    tmp(29042) := x"0062";
    tmp(29043) := x"0062";
    tmp(29044) := x"00a3";
    tmp(29045) := x"00a4";
    tmp(29046) := x"00c4";
    tmp(29047) := x"00c4";
    tmp(29048) := x"08e5";
    tmp(29049) := x"08e5";
    tmp(29050) := x"0905";
    tmp(29051) := x"0905";
    tmp(29052) := x"08e5";
    tmp(29053) := x"0906";
    tmp(29054) := x"08e5";
    tmp(29055) := x"08a4";
    tmp(29056) := x"0082";
    tmp(29057) := x"0042";
    tmp(29058) := x"0021";
    tmp(29059) := x"0020";
    tmp(29060) := x"0020";
    tmp(29061) := x"0020";
    tmp(29062) := x"0020";
    tmp(29063) := x"0041";
    tmp(29064) := x"0883";
    tmp(29065) := x"08a3";
    tmp(29066) := x"00a3";
    tmp(29067) := x"08a3";
    tmp(29068) := x"00a4";
    tmp(29069) := x"08a4";
    tmp(29070) := x"08a4";
    tmp(29071) := x"08a4";
    tmp(29072) := x"08a4";
    tmp(29073) := x"08a3";
    tmp(29074) := x"08c4";
    tmp(29075) := x"08e5";
    tmp(29076) := x"00c4";
    tmp(29077) := x"08c4";
    tmp(29078) := x"08c4";
    tmp(29079) := x"00a3";
    tmp(29080) := x"08e4";
    tmp(29081) := x"08e4";
    tmp(29082) := x"08e4";
    tmp(29083) := x"08e4";
    tmp(29084) := x"08e4";
    tmp(29085) := x"08c4";
    tmp(29086) := x"08a3";
    tmp(29087) := x"08a3";
    tmp(29088) := x"08e4";
    tmp(29089) := x"08e4";
    tmp(29090) := x"0904";
    tmp(29091) := x"0904";
    tmp(29092) := x"08e3";
    tmp(29093) := x"0882";
    tmp(29094) := x"0882";
    tmp(29095) := x"08e4";
    tmp(29096) := x"1125";
    tmp(29097) := x"1166";
    tmp(29098) := x"1125";
    tmp(29099) := x"08c3";
    tmp(29100) := x"10c3";
    tmp(29101) := x"0861";
    tmp(29102) := x"08c2";
    tmp(29103) := x"0905";
    tmp(29104) := x"0987";
    tmp(29105) := x"0967";
    tmp(29106) := x"09c8";
    tmp(29107) := x"124a";
    tmp(29108) := x"124a";
    tmp(29109) := x"1228";
    tmp(29110) := x"1a07";
    tmp(29111) := x"21e6";
    tmp(29112) := x"3a88";
    tmp(29113) := x"636a";
    tmp(29114) := x"83ed";
    tmp(29115) := x"9c6f";
    tmp(29116) := x"acd2";
    tmp(29117) := x"bd74";
    tmp(29118) := x"c5d6";
    tmp(29119) := x"d638";
    tmp(29120) := x"e65a";
    tmp(29121) := x"e69d";
    tmp(29122) := x"e69e";
    tmp(29123) := x"eeff";
    tmp(29124) := x"f71f";
    tmp(29125) := x"f75f";
    tmp(29126) := x"ff9f";
    tmp(29127) := x"ff9f";
    tmp(29128) := x"f79f";
    tmp(29129) := x"ffdf";
    tmp(29130) := x"ffdf";
    tmp(29131) := x"f7df";
    tmp(29132) := x"f7bf";
    tmp(29133) := x"ef9f";
    tmp(29134) := x"ef9f";
    tmp(29135) := x"e79f";
    tmp(29136) := x"e77f";
    tmp(29137) := x"df9f";
    tmp(29138) := x"df7f";
    tmp(29139) := x"cf3f";
    tmp(29140) := x"cf3f";
    tmp(29141) := x"c71f";
    tmp(29142) := x"b69e";
    tmp(29143) := x"ae3c";
    tmp(29144) := x"9d98";
    tmp(29145) := x"9535";
    tmp(29146) := x"9532";
    tmp(29147) := x"7c6e";
    tmp(29148) := x"6bcb";
    tmp(29149) := x"5348";
    tmp(29150) := x"42c5";
    tmp(29151) := x"2a23";
    tmp(29152) := x"19c2";
    tmp(29153) := x"1161";
    tmp(29154) := x"1141";
    tmp(29155) := x"1121";
    tmp(29156) := x"1141";
    tmp(29157) := x"1981";
    tmp(29158) := x"21a2";
    tmp(29159) := x"21c1";
    tmp(29160) := x"19a1";
    tmp(29161) := x"1140";
    tmp(29162) := x"1141";
    tmp(29163) := x"1961";
    tmp(29164) := x"1961";
    tmp(29165) := x"1921";
    tmp(29166) := x"1921";
    tmp(29167) := x"1941";
    tmp(29168) := x"1921";
    tmp(29169) := x"1921";
    tmp(29170) := x"1921";
    tmp(29171) := x"1921";
    tmp(29172) := x"1941";
    tmp(29173) := x"29c1";
    tmp(29174) := x"3a43";
    tmp(29175) := x"52c4";
    tmp(29176) := x"5b26";
    tmp(29177) := x"6346";
    tmp(29178) := x"6b67";
    tmp(29179) := x"7367";
    tmp(29180) := x"7367";
    tmp(29181) := x"7347";
    tmp(29182) := x"6b47";
    tmp(29183) := x"6307";
    tmp(29184) := x"5aa6";
    tmp(29185) := x"4a25";
    tmp(29186) := x"39e3";
    tmp(29187) := x"2982";
    tmp(29188) := x"2141";
    tmp(29189) := x"1921";
    tmp(29190) := x"2121";
    tmp(29191) := x"2141";
    tmp(29192) := x"2141";
    tmp(29193) := x"2141";
    tmp(29194) := x"2961";
    tmp(29195) := x"31a2";
    tmp(29196) := x"3a03";
    tmp(29197) := x"5264";
    tmp(29198) := x"62c6";
    tmp(29199) := x"7b68";
    tmp(29200) := x"8bc9";
    tmp(29201) := x"8bca";
    tmp(29202) := x"83ca";
    tmp(29203) := x"7b89";
    tmp(29204) := x"7348";
    tmp(29205) := x"6b27";
    tmp(29206) := x"62c6";
    tmp(29207) := x"5a86";
    tmp(29208) := x"5a86";
    tmp(29209) := x"5246";
    tmp(29210) := x"4a25";
    tmp(29211) := x"4205";
    tmp(29212) := x"41e5";
    tmp(29213) := x"41c5";
    tmp(29214) := x"41e5";
    tmp(29215) := x"4a26";
    tmp(29216) := x"5267";
    tmp(29217) := x"5a88";
    tmp(29218) := x"62ca";
    tmp(29219) := x"6aeb";
    tmp(29220) := x"7b2d";
    tmp(29221) := x"7b4e";
    tmp(29222) := x"834f";
    tmp(29223) := x"8b70";
    tmp(29224) := x"8bd2";
    tmp(29225) := x"93f4";
    tmp(29226) := x"a435";
    tmp(29227) := x"ac76";
    tmp(29228) := x"ac76";
    tmp(29229) := x"a476";
    tmp(29230) := x"ac76";
    tmp(29231) := x"a456";
    tmp(29232) := x"a476";
    tmp(29233) := x"9c15";
    tmp(29234) := x"a435";
    tmp(29235) := x"a456";
    tmp(29236) := x"9c15";
    tmp(29237) := x"f800";
    tmp(29238) := x"f800";
    tmp(29239) := x"f800";
    tmp(29240) := x"f800";
    tmp(29241) := x"f800";
    tmp(29242) := x"f800";
    tmp(29243) := x"f800";
    tmp(29244) := x"f800";
    tmp(29245) := x"f800";
    tmp(29246) := x"f800";
    tmp(29247) := x"f800";
    tmp(29248) := x"f800";
    tmp(29249) := x"f800";
    tmp(29250) := x"f800";
    tmp(29251) := x"f800";
    tmp(29252) := x"f800";
    tmp(29253) := x"f800";
    tmp(29254) := x"f800";
    tmp(29255) := x"f800";
    tmp(29256) := x"f800";
    tmp(29257) := x"f800";
    tmp(29258) := x"f800";
    tmp(29259) := x"f800";
    tmp(29260) := x"f800";
    tmp(29261) := x"f800";
    tmp(29262) := x"f800";
    tmp(29263) := x"f800";
    tmp(29264) := x"f800";
    tmp(29265) := x"f800";
    tmp(29266) := x"f800";
    tmp(29267) := x"f800";
    tmp(29268) := x"f800";
    tmp(29269) := x"f800";
    tmp(29270) := x"f800";
    tmp(29271) := x"f800";
    tmp(29272) := x"f800";
    tmp(29273) := x"f800";
    tmp(29274) := x"f800";
    tmp(29275) := x"f800";
    tmp(29276) := x"f800";
    tmp(29277) := x"0840";
    tmp(29278) := x"0840";
    tmp(29279) := x"0840";
    tmp(29280) := x"0000";
    tmp(29281) := x"00a4";
    tmp(29282) := x"00c4";
    tmp(29283) := x"00e5";
    tmp(29284) := x"0106";
    tmp(29285) := x"0106";
    tmp(29286) := x"0106";
    tmp(29287) := x"00e5";
    tmp(29288) := x"00e5";
    tmp(29289) := x"00e5";
    tmp(29290) := x"00e5";
    tmp(29291) := x"00e5";
    tmp(29292) := x"00e5";
    tmp(29293) := x"08a4";
    tmp(29294) := x"0041";
    tmp(29295) := x"0021";
    tmp(29296) := x"0020";
    tmp(29297) := x"0000";
    tmp(29298) := x"0020";
    tmp(29299) := x"0020";
    tmp(29300) := x"0020";
    tmp(29301) := x"0020";
    tmp(29302) := x"0041";
    tmp(29303) := x"0862";
    tmp(29304) := x"0882";
    tmp(29305) := x"00a3";
    tmp(29306) := x"08a3";
    tmp(29307) := x"00a3";
    tmp(29308) := x"08a4";
    tmp(29309) := x"08a4";
    tmp(29310) := x"08a4";
    tmp(29311) := x"08a3";
    tmp(29312) := x"08a3";
    tmp(29313) := x"08a3";
    tmp(29314) := x"08e5";
    tmp(29315) := x"08c4";
    tmp(29316) := x"08c4";
    tmp(29317) := x"08c4";
    tmp(29318) := x"08c4";
    tmp(29319) := x"08c4";
    tmp(29320) := x"08c4";
    tmp(29321) := x"0905";
    tmp(29322) := x"08e4";
    tmp(29323) := x"08c4";
    tmp(29324) := x"08c4";
    tmp(29325) := x"08a3";
    tmp(29326) := x"08c4";
    tmp(29327) := x"08c4";
    tmp(29328) := x"0905";
    tmp(29329) := x"0925";
    tmp(29330) := x"08e4";
    tmp(29331) := x"08e4";
    tmp(29332) := x"08e4";
    tmp(29333) := x"08c3";
    tmp(29334) := x"08e4";
    tmp(29335) := x"0904";
    tmp(29336) := x"0905";
    tmp(29337) := x"0925";
    tmp(29338) := x"1145";
    tmp(29339) := x"08c3";
    tmp(29340) := x"08a3";
    tmp(29341) := x"1104";
    tmp(29342) := x"0925";
    tmp(29343) := x"09a8";
    tmp(29344) := x"122a";
    tmp(29345) := x"1229";
    tmp(29346) := x"1207";
    tmp(29347) := x"11a5";
    tmp(29348) := x"1163";
    tmp(29349) := x"1183";
    tmp(29350) := x"21c4";
    tmp(29351) := x"3a25";
    tmp(29352) := x"4a66";
    tmp(29353) := x"5ae7";
    tmp(29354) := x"6b6a";
    tmp(29355) := x"8c0d";
    tmp(29356) := x"944f";
    tmp(29357) := x"acf2";
    tmp(29358) := x"bdb5";
    tmp(29359) := x"c5b7";
    tmp(29360) := x"cdf9";
    tmp(29361) := x"de3b";
    tmp(29362) := x"de5d";
    tmp(29363) := x"e69e";
    tmp(29364) := x"de9f";
    tmp(29365) := x"eedf";
    tmp(29366) := x"f73f";
    tmp(29367) := x"ef1f";
    tmp(29368) := x"ef3f";
    tmp(29369) := x"ef5f";
    tmp(29370) := x"ef7f";
    tmp(29371) := x"df1f";
    tmp(29372) := x"e71f";
    tmp(29373) := x"df1f";
    tmp(29374) := x"df3f";
    tmp(29375) := x"df1f";
    tmp(29376) := x"d6ff";
    tmp(29377) := x"d71f";
    tmp(29378) := x"d73f";
    tmp(29379) := x"cf1f";
    tmp(29380) := x"be9f";
    tmp(29381) := x"b63d";
    tmp(29382) := x"adfb";
    tmp(29383) := x"9dd9";
    tmp(29384) := x"9534";
    tmp(29385) := x"8cd2";
    tmp(29386) := x"848f";
    tmp(29387) := x"6beb";
    tmp(29388) := x"5b69";
    tmp(29389) := x"42c6";
    tmp(29390) := x"3244";
    tmp(29391) := x"21a2";
    tmp(29392) := x"1182";
    tmp(29393) := x"1161";
    tmp(29394) := x"1141";
    tmp(29395) := x"1141";
    tmp(29396) := x"1962";
    tmp(29397) := x"19a2";
    tmp(29398) := x"21c2";
    tmp(29399) := x"21c1";
    tmp(29400) := x"1961";
    tmp(29401) := x"1140";
    tmp(29402) := x"1140";
    tmp(29403) := x"1141";
    tmp(29404) := x"1961";
    tmp(29405) := x"1941";
    tmp(29406) := x"1941";
    tmp(29407) := x"1941";
    tmp(29408) := x"1941";
    tmp(29409) := x"1942";
    tmp(29410) := x"1942";
    tmp(29411) := x"1921";
    tmp(29412) := x"1921";
    tmp(29413) := x"1961";
    tmp(29414) := x"29e1";
    tmp(29415) := x"4263";
    tmp(29416) := x"52c4";
    tmp(29417) := x"5ae5";
    tmp(29418) := x"6326";
    tmp(29419) := x"6b26";
    tmp(29420) := x"6b47";
    tmp(29421) := x"6b47";
    tmp(29422) := x"6b47";
    tmp(29423) := x"6b27";
    tmp(29424) := x"62e6";
    tmp(29425) := x"5285";
    tmp(29426) := x"4224";
    tmp(29427) := x"39e3";
    tmp(29428) := x"2982";
    tmp(29429) := x"2121";
    tmp(29430) := x"1901";
    tmp(29431) := x"2121";
    tmp(29432) := x"2141";
    tmp(29433) := x"2141";
    tmp(29434) := x"2161";
    tmp(29435) := x"2961";
    tmp(29436) := x"31a2";
    tmp(29437) := x"39e3";
    tmp(29438) := x"4a44";
    tmp(29439) := x"5aa6";
    tmp(29440) := x"7b48";
    tmp(29441) := x"8389";
    tmp(29442) := x"7b68";
    tmp(29443) := x"7368";
    tmp(29444) := x"6b28";
    tmp(29445) := x"6ae7";
    tmp(29446) := x"5aa6";
    tmp(29447) := x"5265";
    tmp(29448) := x"5245";
    tmp(29449) := x"4a05";
    tmp(29450) := x"41e4";
    tmp(29451) := x"39a4";
    tmp(29452) := x"39a4";
    tmp(29453) := x"39a4";
    tmp(29454) := x"41e5";
    tmp(29455) := x"4a06";
    tmp(29456) := x"5247";
    tmp(29457) := x"5a68";
    tmp(29458) := x"5a89";
    tmp(29459) := x"628a";
    tmp(29460) := x"72cb";
    tmp(29461) := x"730c";
    tmp(29462) := x"7b2d";
    tmp(29463) := x"834f";
    tmp(29464) := x"8b90";
    tmp(29465) := x"93d2";
    tmp(29466) := x"93f3";
    tmp(29467) := x"a434";
    tmp(29468) := x"a456";
    tmp(29469) := x"a456";
    tmp(29470) := x"a456";
    tmp(29471) := x"a456";
    tmp(29472) := x"a476";
    tmp(29473) := x"9c35";
    tmp(29474) := x"a435";
    tmp(29475) := x"a435";
    tmp(29476) := x"9bf5";
    tmp(29477) := x"f800";
    tmp(29478) := x"f800";
    tmp(29479) := x"f800";
    tmp(29480) := x"f800";
    tmp(29481) := x"f800";
    tmp(29482) := x"f800";
    tmp(29483) := x"f800";
    tmp(29484) := x"f800";
    tmp(29485) := x"f800";
    tmp(29486) := x"f800";
    tmp(29487) := x"f800";
    tmp(29488) := x"f800";
    tmp(29489) := x"f800";
    tmp(29490) := x"f800";
    tmp(29491) := x"f800";
    tmp(29492) := x"f800";
    tmp(29493) := x"f800";
    tmp(29494) := x"f800";
    tmp(29495) := x"f800";
    tmp(29496) := x"f800";
    tmp(29497) := x"f800";
    tmp(29498) := x"f800";
    tmp(29499) := x"f800";
    tmp(29500) := x"f800";
    tmp(29501) := x"f800";
    tmp(29502) := x"f800";
    tmp(29503) := x"f800";
    tmp(29504) := x"f800";
    tmp(29505) := x"f800";
    tmp(29506) := x"f800";
    tmp(29507) := x"f800";
    tmp(29508) := x"f800";
    tmp(29509) := x"f800";
    tmp(29510) := x"f800";
    tmp(29511) := x"f800";
    tmp(29512) := x"f800";
    tmp(29513) := x"f800";
    tmp(29514) := x"f800";
    tmp(29515) := x"f800";
    tmp(29516) := x"f800";
    tmp(29517) := x"0840";
    tmp(29518) := x"0840";
    tmp(29519) := x"0840";
    tmp(29520) := x"0020";
    tmp(29521) := x"00e5";
    tmp(29522) := x"00e5";
    tmp(29523) := x"00e5";
    tmp(29524) := x"00e5";
    tmp(29525) := x"00e5";
    tmp(29526) := x"00e5";
    tmp(29527) := x"00c5";
    tmp(29528) := x"00c5";
    tmp(29529) := x"00c5";
    tmp(29530) := x"00e5";
    tmp(29531) := x"00e5";
    tmp(29532) := x"00a4";
    tmp(29533) := x"0021";
    tmp(29534) := x"0020";
    tmp(29535) := x"0000";
    tmp(29536) := x"0020";
    tmp(29537) := x"0020";
    tmp(29538) := x"0021";
    tmp(29539) := x"0841";
    tmp(29540) := x"0021";
    tmp(29541) := x"0861";
    tmp(29542) := x"0882";
    tmp(29543) := x"08a3";
    tmp(29544) := x"0883";
    tmp(29545) := x"08a4";
    tmp(29546) := x"08a4";
    tmp(29547) := x"08c4";
    tmp(29548) := x"08c4";
    tmp(29549) := x"08c4";
    tmp(29550) := x"08a4";
    tmp(29551) := x"08a4";
    tmp(29552) := x"08a4";
    tmp(29553) := x"08e4";
    tmp(29554) := x"08e5";
    tmp(29555) := x"08e5";
    tmp(29556) := x"08c4";
    tmp(29557) := x"08c4";
    tmp(29558) := x"08e4";
    tmp(29559) := x"08e4";
    tmp(29560) := x"08e4";
    tmp(29561) := x"08e4";
    tmp(29562) := x"08e4";
    tmp(29563) := x"08c3";
    tmp(29564) := x"08c4";
    tmp(29565) := x"08c4";
    tmp(29566) := x"08e4";
    tmp(29567) := x"08c4";
    tmp(29568) := x"08e4";
    tmp(29569) := x"0925";
    tmp(29570) := x"0905";
    tmp(29571) := x"08c3";
    tmp(29572) := x"08c3";
    tmp(29573) := x"08c3";
    tmp(29574) := x"08c3";
    tmp(29575) := x"08e4";
    tmp(29576) := x"0904";
    tmp(29577) := x"0925";
    tmp(29578) := x"1146";
    tmp(29579) := x"1104";
    tmp(29580) := x"1105";
    tmp(29581) := x"19c7";
    tmp(29582) := x"11a6";
    tmp(29583) := x"09c6";
    tmp(29584) := x"09a5";
    tmp(29585) := x"0963";
    tmp(29586) := x"0921";
    tmp(29587) := x"0901";
    tmp(29588) := x"1101";
    tmp(29589) := x"1941";
    tmp(29590) := x"2182";
    tmp(29591) := x"31e4";
    tmp(29592) := x"3a45";
    tmp(29593) := x"4a86";
    tmp(29594) := x"6308";
    tmp(29595) := x"736b";
    tmp(29596) := x"8bee";
    tmp(29597) := x"a491";
    tmp(29598) := x"acf2";
    tmp(29599) := x"bd76";
    tmp(29600) := x"c5b8";
    tmp(29601) := x"c5b9";
    tmp(29602) := x"cddb";
    tmp(29603) := x"cddc";
    tmp(29604) := x"d61e";
    tmp(29605) := x"de9f";
    tmp(29606) := x"de9f";
    tmp(29607) := x"de9f";
    tmp(29608) := x"de9f";
    tmp(29609) := x"debf";
    tmp(29610) := x"e71f";
    tmp(29611) := x"d69f";
    tmp(29612) := x"ce9f";
    tmp(29613) := x"ce5f";
    tmp(29614) := x"d69f";
    tmp(29615) := x"c67f";
    tmp(29616) := x"c65f";
    tmp(29617) := x"c69f";
    tmp(29618) := x"c69f";
    tmp(29619) := x"be7e";
    tmp(29620) := x"ae1d";
    tmp(29621) := x"a5da";
    tmp(29622) := x"a598";
    tmp(29623) := x"9535";
    tmp(29624) := x"8cd2";
    tmp(29625) := x"846f";
    tmp(29626) := x"73ec";
    tmp(29627) := x"5b49";
    tmp(29628) := x"4ac6";
    tmp(29629) := x"3a85";
    tmp(29630) := x"21e3";
    tmp(29631) := x"1982";
    tmp(29632) := x"1162";
    tmp(29633) := x"1162";
    tmp(29634) := x"1162";
    tmp(29635) := x"1982";
    tmp(29636) := x"19a2";
    tmp(29637) := x"21c2";
    tmp(29638) := x"29e2";
    tmp(29639) := x"19a1";
    tmp(29640) := x"1120";
    tmp(29641) := x"1120";
    tmp(29642) := x"1140";
    tmp(29643) := x"1141";
    tmp(29644) := x"1961";
    tmp(29645) := x"1961";
    tmp(29646) := x"1941";
    tmp(29647) := x"1941";
    tmp(29648) := x"1942";
    tmp(29649) := x"1962";
    tmp(29650) := x"1942";
    tmp(29651) := x"1941";
    tmp(29652) := x"1921";
    tmp(29653) := x"1921";
    tmp(29654) := x"2181";
    tmp(29655) := x"3202";
    tmp(29656) := x"4263";
    tmp(29657) := x"52c4";
    tmp(29658) := x"5ae5";
    tmp(29659) := x"6306";
    tmp(29660) := x"6306";
    tmp(29661) := x"6b26";
    tmp(29662) := x"6b26";
    tmp(29663) := x"6306";
    tmp(29664) := x"62e6";
    tmp(29665) := x"5ac6";
    tmp(29666) := x"5265";
    tmp(29667) := x"4224";
    tmp(29668) := x"31c3";
    tmp(29669) := x"2962";
    tmp(29670) := x"2121";
    tmp(29671) := x"2121";
    tmp(29672) := x"2121";
    tmp(29673) := x"2141";
    tmp(29674) := x"2141";
    tmp(29675) := x"2961";
    tmp(29676) := x"2982";
    tmp(29677) := x"3182";
    tmp(29678) := x"39e3";
    tmp(29679) := x"4a24";
    tmp(29680) := x"62a6";
    tmp(29681) := x"6b07";
    tmp(29682) := x"7328";
    tmp(29683) := x"6b28";
    tmp(29684) := x"6ae7";
    tmp(29685) := x"5aa6";
    tmp(29686) := x"5285";
    tmp(29687) := x"4a25";
    tmp(29688) := x"41e4";
    tmp(29689) := x"41e4";
    tmp(29690) := x"39a4";
    tmp(29691) := x"3183";
    tmp(29692) := x"3184";
    tmp(29693) := x"3984";
    tmp(29694) := x"39c5";
    tmp(29695) := x"41e6";
    tmp(29696) := x"49e6";
    tmp(29697) := x"5207";
    tmp(29698) := x"5248";
    tmp(29699) := x"5a69";
    tmp(29700) := x"6aaa";
    tmp(29701) := x"6acb";
    tmp(29702) := x"6acd";
    tmp(29703) := x"7b0e";
    tmp(29704) := x"834f";
    tmp(29705) := x"8b91";
    tmp(29706) := x"8bb2";
    tmp(29707) := x"93f3";
    tmp(29708) := x"a475";
    tmp(29709) := x"a456";
    tmp(29710) := x"ac76";
    tmp(29711) := x"a456";
    tmp(29712) := x"ac76";
    tmp(29713) := x"a455";
    tmp(29714) := x"9c15";
    tmp(29715) := x"a456";
    tmp(29716) := x"a415";
    tmp(29717) := x"f800";
    tmp(29718) := x"f800";
    tmp(29719) := x"f800";
    tmp(29720) := x"f800";
    tmp(29721) := x"f800";
    tmp(29722) := x"f800";
    tmp(29723) := x"f800";
    tmp(29724) := x"f800";
    tmp(29725) := x"f800";
    tmp(29726) := x"f800";
    tmp(29727) := x"f800";
    tmp(29728) := x"f800";
    tmp(29729) := x"f800";
    tmp(29730) := x"f800";
    tmp(29731) := x"f800";
    tmp(29732) := x"f800";
    tmp(29733) := x"f800";
    tmp(29734) := x"f800";
    tmp(29735) := x"f800";
    tmp(29736) := x"f800";
    tmp(29737) := x"f800";
    tmp(29738) := x"f800";
    tmp(29739) := x"f800";
    tmp(29740) := x"f800";
    tmp(29741) := x"f800";
    tmp(29742) := x"f800";
    tmp(29743) := x"f800";
    tmp(29744) := x"f800";
    tmp(29745) := x"f800";
    tmp(29746) := x"f800";
    tmp(29747) := x"f800";
    tmp(29748) := x"f800";
    tmp(29749) := x"f800";
    tmp(29750) := x"f800";
    tmp(29751) := x"f800";
    tmp(29752) := x"f800";
    tmp(29753) := x"f800";
    tmp(29754) := x"f800";
    tmp(29755) := x"f800";
    tmp(29756) := x"f800";
    tmp(29757) := x"0840";
    tmp(29758) := x"0840";
    tmp(29759) := x"0840";
    tmp(29760) := x"0020";
    tmp(29761) := x"00c5";
    tmp(29762) := x"00c5";
    tmp(29763) := x"00c5";
    tmp(29764) := x"00c5";
    tmp(29765) := x"00e5";
    tmp(29766) := x"00e5";
    tmp(29767) := x"00e5";
    tmp(29768) := x"00c5";
    tmp(29769) := x"00e5";
    tmp(29770) := x"00e5";
    tmp(29771) := x"00e5";
    tmp(29772) := x"00a4";
    tmp(29773) := x"0041";
    tmp(29774) := x"0020";
    tmp(29775) := x"0020";
    tmp(29776) := x"0020";
    tmp(29777) := x"0021";
    tmp(29778) := x"0062";
    tmp(29779) := x"0882";
    tmp(29780) := x"0862";
    tmp(29781) := x"08a3";
    tmp(29782) := x"08c4";
    tmp(29783) := x"08c4";
    tmp(29784) := x"08a4";
    tmp(29785) := x"08c4";
    tmp(29786) := x"08a4";
    tmp(29787) := x"08c5";
    tmp(29788) := x"08e5";
    tmp(29789) := x"08e5";
    tmp(29790) := x"08e5";
    tmp(29791) := x"08c4";
    tmp(29792) := x"08c4";
    tmp(29793) := x"08e5";
    tmp(29794) := x"0905";
    tmp(29795) := x"0905";
    tmp(29796) := x"08e4";
    tmp(29797) := x"08e4";
    tmp(29798) := x"08e4";
    tmp(29799) := x"0905";
    tmp(29800) := x"08e4";
    tmp(29801) := x"08e4";
    tmp(29802) := x"08e4";
    tmp(29803) := x"08c3";
    tmp(29804) := x"08e4";
    tmp(29805) := x"08e4";
    tmp(29806) := x"08e4";
    tmp(29807) := x"08c3";
    tmp(29808) := x"08c3";
    tmp(29809) := x"08c4";
    tmp(29810) := x"0905";
    tmp(29811) := x"08e4";
    tmp(29812) := x"08c3";
    tmp(29813) := x"08c3";
    tmp(29814) := x"08e4";
    tmp(29815) := x"0904";
    tmp(29816) := x"0904";
    tmp(29817) := x"0904";
    tmp(29818) := x"1145";
    tmp(29819) := x"0882";
    tmp(29820) := x"08e4";
    tmp(29821) := x"11c6";
    tmp(29822) := x"0902";
    tmp(29823) := x"0901";
    tmp(29824) := x"08c0";
    tmp(29825) := x"08c0";
    tmp(29826) := x"08c0";
    tmp(29827) := x"08e0";
    tmp(29828) := x"1101";
    tmp(29829) := x"1121";
    tmp(29830) := x"1962";
    tmp(29831) := x"29a3";
    tmp(29832) := x"3a04";
    tmp(29833) := x"4245";
    tmp(29834) := x"52a7";
    tmp(29835) := x"6309";
    tmp(29836) := x"7b8c";
    tmp(29837) := x"8c0f";
    tmp(29838) := x"9c91";
    tmp(29839) := x"acf3";
    tmp(29840) := x"b536";
    tmp(29841) := x"bd78";
    tmp(29842) := x"bd79";
    tmp(29843) := x"c59a";
    tmp(29844) := x"c5bc";
    tmp(29845) := x"cdfc";
    tmp(29846) := x"ce1e";
    tmp(29847) := x"c5fe";
    tmp(29848) := x"c63f";
    tmp(29849) := x"c63e";
    tmp(29850) := x"ce5e";
    tmp(29851) := x"c63f";
    tmp(29852) := x"c61f";
    tmp(29853) := x"bdff";
    tmp(29854) := x"c63f";
    tmp(29855) := x"be3f";
    tmp(29856) := x"be3f";
    tmp(29857) := x"b61f";
    tmp(29858) := x"b5fe";
    tmp(29859) := x"addd";
    tmp(29860) := x"a5bb";
    tmp(29861) := x"9d57";
    tmp(29862) := x"9515";
    tmp(29863) := x"8cb2";
    tmp(29864) := x"846f";
    tmp(29865) := x"73ec";
    tmp(29866) := x"636a";
    tmp(29867) := x"52c7";
    tmp(29868) := x"3a65";
    tmp(29869) := x"2a03";
    tmp(29870) := x"1982";
    tmp(29871) := x"1162";
    tmp(29872) := x"1142";
    tmp(29873) := x"1162";
    tmp(29874) := x"1982";
    tmp(29875) := x"19a2";
    tmp(29876) := x"21c3";
    tmp(29877) := x"29e3";
    tmp(29878) := x"2a02";
    tmp(29879) := x"1961";
    tmp(29880) := x"1120";
    tmp(29881) := x"1120";
    tmp(29882) := x"1120";
    tmp(29883) := x"1140";
    tmp(29884) := x"1141";
    tmp(29885) := x"1961";
    tmp(29886) := x"1961";
    tmp(29887) := x"1961";
    tmp(29888) := x"1962";
    tmp(29889) := x"1962";
    tmp(29890) := x"1962";
    tmp(29891) := x"1942";
    tmp(29892) := x"1921";
    tmp(29893) := x"1101";
    tmp(29894) := x"1921";
    tmp(29895) := x"2181";
    tmp(29896) := x"3202";
    tmp(29897) := x"4263";
    tmp(29898) := x"52a4";
    tmp(29899) := x"52c5";
    tmp(29900) := x"5ae5";
    tmp(29901) := x"62e6";
    tmp(29902) := x"6306";
    tmp(29903) := x"6306";
    tmp(29904) := x"5ac6";
    tmp(29905) := x"5ac6";
    tmp(29906) := x"5aa5";
    tmp(29907) := x"4a45";
    tmp(29908) := x"4204";
    tmp(29909) := x"31a3";
    tmp(29910) := x"2942";
    tmp(29911) := x"2121";
    tmp(29912) := x"2121";
    tmp(29913) := x"2141";
    tmp(29914) := x"2141";
    tmp(29915) := x"2961";
    tmp(29916) := x"2962";
    tmp(29917) := x"2982";
    tmp(29918) := x"3182";
    tmp(29919) := x"39e3";
    tmp(29920) := x"4a44";
    tmp(29921) := x"62a6";
    tmp(29922) := x"6ac7";
    tmp(29923) := x"6ac7";
    tmp(29924) := x"62a6";
    tmp(29925) := x"5285";
    tmp(29926) := x"4a45";
    tmp(29927) := x"41e4";
    tmp(29928) := x"39c3";
    tmp(29929) := x"39a4";
    tmp(29930) := x"3163";
    tmp(29931) := x"3163";
    tmp(29932) := x"3163";
    tmp(29933) := x"3184";
    tmp(29934) := x"39a5";
    tmp(29935) := x"39a5";
    tmp(29936) := x"41c6";
    tmp(29937) := x"41c6";
    tmp(29938) := x"5207";
    tmp(29939) := x"5248";
    tmp(29940) := x"5a69";
    tmp(29941) := x"628a";
    tmp(29942) := x"6a8c";
    tmp(29943) := x"6acd";
    tmp(29944) := x"730e";
    tmp(29945) := x"834f";
    tmp(29946) := x"8371";
    tmp(29947) := x"8bd2";
    tmp(29948) := x"93f3";
    tmp(29949) := x"9c15";
    tmp(29950) := x"a435";
    tmp(29951) := x"a476";
    tmp(29952) := x"ac77";
    tmp(29953) := x"a436";
    tmp(29954) := x"9c36";
    tmp(29955) := x"9c35";
    tmp(29956) := x"93d4";
    tmp(29957) := x"07e0";
    tmp(29958) := x"07e0";
    tmp(29959) := x"07e0";
    tmp(29960) := x"07e0";
    tmp(29961) := x"07e0";
    tmp(29962) := x"07e0";
    tmp(29963) := x"07e0";
    tmp(29964) := x"07e0";
    tmp(29965) := x"07e0";
    tmp(29966) := x"07e0";
    tmp(29967) := x"07e0";
    tmp(29968) := x"07e0";
    tmp(29969) := x"07e0";
    tmp(29970) := x"07e0";
    tmp(29971) := x"07e0";
    tmp(29972) := x"07e0";
    tmp(29973) := x"07e0";
    tmp(29974) := x"07e0";
    tmp(29975) := x"07e0";
    tmp(29976) := x"07e0";
    tmp(29977) := x"07e0";
    tmp(29978) := x"07e0";
    tmp(29979) := x"07e0";
    tmp(29980) := x"07e0";
    tmp(29981) := x"07e0";
    tmp(29982) := x"07e0";
    tmp(29983) := x"07e0";
    tmp(29984) := x"07e0";
    tmp(29985) := x"07e0";
    tmp(29986) := x"07e0";
    tmp(29987) := x"07e0";
    tmp(29988) := x"07e0";
    tmp(29989) := x"07e0";
    tmp(29990) := x"07e0";
    tmp(29991) := x"07e0";
    tmp(29992) := x"07e0";
    tmp(29993) := x"07e0";
    tmp(29994) := x"07e0";
    tmp(29995) := x"07e0";
    tmp(29996) := x"07e0";
    tmp(29997) := x"0840";
    tmp(29998) := x"0840";
    tmp(29999) := x"0840";
    tmp(30000) := x"0020";
    tmp(30001) := x"00c5";
    tmp(30002) := x"00c5";
    tmp(30003) := x"00e5";
    tmp(30004) := x"00c5";
    tmp(30005) := x"00e5";
    tmp(30006) := x"00e5";
    tmp(30007) := x"00e5";
    tmp(30008) := x"00e5";
    tmp(30009) := x"00e5";
    tmp(30010) := x"00e5";
    tmp(30011) := x"00a3";
    tmp(30012) := x"0041";
    tmp(30013) := x"0021";
    tmp(30014) := x"0021";
    tmp(30015) := x"0841";
    tmp(30016) := x"0861";
    tmp(30017) := x"0882";
    tmp(30018) := x"08c4";
    tmp(30019) := x"08e5";
    tmp(30020) := x"08e5";
    tmp(30021) := x"0905";
    tmp(30022) := x"0906";
    tmp(30023) := x"0906";
    tmp(30024) := x"0906";
    tmp(30025) := x"0906";
    tmp(30026) := x"0906";
    tmp(30027) := x"08e5";
    tmp(30028) := x"08c5";
    tmp(30029) := x"08c5";
    tmp(30030) := x"08c5";
    tmp(30031) := x"08c5";
    tmp(30032) := x"08c5";
    tmp(30033) := x"08e5";
    tmp(30034) := x"08c4";
    tmp(30035) := x"08e4";
    tmp(30036) := x"08e4";
    tmp(30037) := x"08e4";
    tmp(30038) := x"08c4";
    tmp(30039) := x"08e5";
    tmp(30040) := x"0905";
    tmp(30041) := x"0905";
    tmp(30042) := x"08e4";
    tmp(30043) := x"08e4";
    tmp(30044) := x"0904";
    tmp(30045) := x"08e4";
    tmp(30046) := x"08e4";
    tmp(30047) := x"08e4";
    tmp(30048) := x"08a3";
    tmp(30049) := x"0883";
    tmp(30050) := x"08e4";
    tmp(30051) := x"08e4";
    tmp(30052) := x"08e4";
    tmp(30053) := x"08e3";
    tmp(30054) := x"0904";
    tmp(30055) := x"0904";
    tmp(30056) := x"0904";
    tmp(30057) := x"0904";
    tmp(30058) := x"08e4";
    tmp(30059) := x"0882";
    tmp(30060) := x"0904";
    tmp(30061) := x"19c6";
    tmp(30062) := x"08c1";
    tmp(30063) := x"08a0";
    tmp(30064) := x"08c0";
    tmp(30065) := x"08c0";
    tmp(30066) := x"08c0";
    tmp(30067) := x"08c0";
    tmp(30068) := x"0900";
    tmp(30069) := x"1101";
    tmp(30070) := x"1941";
    tmp(30071) := x"2182";
    tmp(30072) := x"29c3";
    tmp(30073) := x"3a25";
    tmp(30074) := x"4246";
    tmp(30075) := x"52a8";
    tmp(30076) := x"630a";
    tmp(30077) := x"7bad";
    tmp(30078) := x"8c0e";
    tmp(30079) := x"9c91";
    tmp(30080) := x"a4d3";
    tmp(30081) := x"acf5";
    tmp(30082) := x"b517";
    tmp(30083) := x"b538";
    tmp(30084) := x"bd7a";
    tmp(30085) := x"bd9b";
    tmp(30086) := x"bd9c";
    tmp(30087) := x"bdbd";
    tmp(30088) := x"bdfc";
    tmp(30089) := x"b5bc";
    tmp(30090) := x"bddd";
    tmp(30091) := x"b59c";
    tmp(30092) := x"b5bd";
    tmp(30093) := x"b5bd";
    tmp(30094) := x"b5be";
    tmp(30095) := x"b5bd";
    tmp(30096) := x"adbd";
    tmp(30097) := x"a5bd";
    tmp(30098) := x"a57b";
    tmp(30099) := x"9d59";
    tmp(30100) := x"9517";
    tmp(30101) := x"8cd4";
    tmp(30102) := x"8cb2";
    tmp(30103) := x"742e";
    tmp(30104) := x"6bcc";
    tmp(30105) := x"634a";
    tmp(30106) := x"52e7";
    tmp(30107) := x"3a65";
    tmp(30108) := x"2a04";
    tmp(30109) := x"19a3";
    tmp(30110) := x"1162";
    tmp(30111) := x"1162";
    tmp(30112) := x"1162";
    tmp(30113) := x"1182";
    tmp(30114) := x"19a3";
    tmp(30115) := x"21c3";
    tmp(30116) := x"2a03";
    tmp(30117) := x"2a23";
    tmp(30118) := x"21c1";
    tmp(30119) := x"1141";
    tmp(30120) := x"1120";
    tmp(30121) := x"1120";
    tmp(30122) := x"1120";
    tmp(30123) := x"1120";
    tmp(30124) := x"1141";
    tmp(30125) := x"1941";
    tmp(30126) := x"1961";
    tmp(30127) := x"1961";
    tmp(30128) := x"1962";
    tmp(30129) := x"1983";
    tmp(30130) := x"1963";
    tmp(30131) := x"1962";
    tmp(30132) := x"1941";
    tmp(30133) := x"1121";
    tmp(30134) := x"1921";
    tmp(30135) := x"1941";
    tmp(30136) := x"21a1";
    tmp(30137) := x"3202";
    tmp(30138) := x"4263";
    tmp(30139) := x"4a84";
    tmp(30140) := x"52a4";
    tmp(30141) := x"5ac5";
    tmp(30142) := x"5ac5";
    tmp(30143) := x"5ac5";
    tmp(30144) := x"5aa5";
    tmp(30145) := x"5aa5";
    tmp(30146) := x"5aa5";
    tmp(30147) := x"5265";
    tmp(30148) := x"4a45";
    tmp(30149) := x"39e4";
    tmp(30150) := x"3182";
    tmp(30151) := x"2142";
    tmp(30152) := x"2121";
    tmp(30153) := x"2121";
    tmp(30154) := x"2141";
    tmp(30155) := x"2161";
    tmp(30156) := x"2962";
    tmp(30157) := x"2962";
    tmp(30158) := x"2982";
    tmp(30159) := x"31a2";
    tmp(30160) := x"39c3";
    tmp(30161) := x"4a24";
    tmp(30162) := x"5a86";
    tmp(30163) := x"5a86";
    tmp(30164) := x"5266";
    tmp(30165) := x"5245";
    tmp(30166) := x"4a24";
    tmp(30167) := x"41e4";
    tmp(30168) := x"3183";
    tmp(30169) := x"3163";
    tmp(30170) := x"2943";
    tmp(30171) := x"2943";
    tmp(30172) := x"2943";
    tmp(30173) := x"3163";
    tmp(30174) := x"3184";
    tmp(30175) := x"3984";
    tmp(30176) := x"39a5";
    tmp(30177) := x"41c6";
    tmp(30178) := x"41e6";
    tmp(30179) := x"5207";
    tmp(30180) := x"5228";
    tmp(30181) := x"5a49";
    tmp(30182) := x"5a4a";
    tmp(30183) := x"6a8b";
    tmp(30184) := x"72cd";
    tmp(30185) := x"730d";
    tmp(30186) := x"7b4f";
    tmp(30187) := x"8b91";
    tmp(30188) := x"93d2";
    tmp(30189) := x"9bf3";
    tmp(30190) := x"9c34";
    tmp(30191) := x"9c55";
    tmp(30192) := x"a456";
    tmp(30193) := x"9c15";
    tmp(30194) := x"9c14";
    tmp(30195) := x"9c15";
    tmp(30196) := x"93d4";
    tmp(30197) := x"07e0";
    tmp(30198) := x"07e0";
    tmp(30199) := x"07e0";
    tmp(30200) := x"07e0";
    tmp(30201) := x"07e0";
    tmp(30202) := x"07e0";
    tmp(30203) := x"07e0";
    tmp(30204) := x"07e0";
    tmp(30205) := x"07e0";
    tmp(30206) := x"07e0";
    tmp(30207) := x"07e0";
    tmp(30208) := x"07e0";
    tmp(30209) := x"07e0";
    tmp(30210) := x"07e0";
    tmp(30211) := x"07e0";
    tmp(30212) := x"07e0";
    tmp(30213) := x"07e0";
    tmp(30214) := x"07e0";
    tmp(30215) := x"07e0";
    tmp(30216) := x"07e0";
    tmp(30217) := x"07e0";
    tmp(30218) := x"07e0";
    tmp(30219) := x"07e0";
    tmp(30220) := x"07e0";
    tmp(30221) := x"07e0";
    tmp(30222) := x"07e0";
    tmp(30223) := x"07e0";
    tmp(30224) := x"07e0";
    tmp(30225) := x"07e0";
    tmp(30226) := x"07e0";
    tmp(30227) := x"07e0";
    tmp(30228) := x"07e0";
    tmp(30229) := x"07e0";
    tmp(30230) := x"07e0";
    tmp(30231) := x"07e0";
    tmp(30232) := x"07e0";
    tmp(30233) := x"07e0";
    tmp(30234) := x"07e0";
    tmp(30235) := x"07e0";
    tmp(30236) := x"07e0";
    tmp(30237) := x"0840";
    tmp(30238) := x"0840";
    tmp(30239) := x"0840";
    tmp(30240) := x"0000";
    tmp(30241) := x"00c4";
    tmp(30242) := x"00a4";
    tmp(30243) := x"00c4";
    tmp(30244) := x"00c4";
    tmp(30245) := x"00e5";
    tmp(30246) := x"00e5";
    tmp(30247) := x"00e6";
    tmp(30248) := x"0106";
    tmp(30249) := x"0106";
    tmp(30250) := x"08e6";
    tmp(30251) := x"0041";
    tmp(30252) := x"0020";
    tmp(30253) := x"0020";
    tmp(30254) := x"0021";
    tmp(30255) := x"0862";
    tmp(30256) := x"08a3";
    tmp(30257) := x"08c4";
    tmp(30258) := x"08c4";
    tmp(30259) := x"08e5";
    tmp(30260) := x"08e5";
    tmp(30261) := x"08e5";
    tmp(30262) := x"08c5";
    tmp(30263) := x"08c5";
    tmp(30264) := x"08a4";
    tmp(30265) := x"08a4";
    tmp(30266) := x"08a3";
    tmp(30267) := x"08a3";
    tmp(30268) := x"08a3";
    tmp(30269) := x"0883";
    tmp(30270) := x"08a4";
    tmp(30271) := x"08a4";
    tmp(30272) := x"08c4";
    tmp(30273) := x"08c4";
    tmp(30274) := x"08c4";
    tmp(30275) := x"08c4";
    tmp(30276) := x"08e4";
    tmp(30277) := x"08c4";
    tmp(30278) := x"08e5";
    tmp(30279) := x"08e5";
    tmp(30280) := x"08e5";
    tmp(30281) := x"0905";
    tmp(30282) := x"0905";
    tmp(30283) := x"0905";
    tmp(30284) := x"0926";
    tmp(30285) := x"0905";
    tmp(30286) := x"0905";
    tmp(30287) := x"0882";
    tmp(30288) := x"0862";
    tmp(30289) := x"08a3";
    tmp(30290) := x"08e4";
    tmp(30291) := x"08e4";
    tmp(30292) := x"0904";
    tmp(30293) := x"0904";
    tmp(30294) := x"08e4";
    tmp(30295) := x"0925";
    tmp(30296) := x"0904";
    tmp(30297) := x"0904";
    tmp(30298) := x"08a3";
    tmp(30299) := x"08a3";
    tmp(30300) := x"1125";
    tmp(30301) := x"19c5";
    tmp(30302) := x"08a0";
    tmp(30303) := x"08c0";
    tmp(30304) := x"08c0";
    tmp(30305) := x"08c0";
    tmp(30306) := x"08c0";
    tmp(30307) := x"08c0";
    tmp(30308) := x"08e0";
    tmp(30309) := x"08e1";
    tmp(30310) := x"1121";
    tmp(30311) := x"1962";
    tmp(30312) := x"21a2";
    tmp(30313) := x"31e4";
    tmp(30314) := x"3a25";
    tmp(30315) := x"4246";
    tmp(30316) := x"52c9";
    tmp(30317) := x"6b4b";
    tmp(30318) := x"7bad";
    tmp(30319) := x"8c0f";
    tmp(30320) := x"9471";
    tmp(30321) := x"a4b3";
    tmp(30322) := x"a4b4";
    tmp(30323) := x"a4d6";
    tmp(30324) := x"a4f7";
    tmp(30325) := x"b539";
    tmp(30326) := x"ad39";
    tmp(30327) := x"b53a";
    tmp(30328) := x"ad7a";
    tmp(30329) := x"ad7b";
    tmp(30330) := x"ad1a";
    tmp(30331) := x"a53b";
    tmp(30332) := x"a51a";
    tmp(30333) := x"a53b";
    tmp(30334) := x"a57c";
    tmp(30335) := x"a55c";
    tmp(30336) := x"9d5b";
    tmp(30337) := x"9d3a";
    tmp(30338) := x"94f8";
    tmp(30339) := x"8cd5";
    tmp(30340) := x"8473";
    tmp(30341) := x"7c31";
    tmp(30342) := x"7c0e";
    tmp(30343) := x"6bac";
    tmp(30344) := x"6349";
    tmp(30345) := x"5307";
    tmp(30346) := x"4265";
    tmp(30347) := x"3204";
    tmp(30348) := x"21a3";
    tmp(30349) := x"1962";
    tmp(30350) := x"1162";
    tmp(30351) := x"1162";
    tmp(30352) := x"1183";
    tmp(30353) := x"19a3";
    tmp(30354) := x"21a3";
    tmp(30355) := x"2a03";
    tmp(30356) := x"3244";
    tmp(30357) := x"2a23";
    tmp(30358) := x"1981";
    tmp(30359) := x"1120";
    tmp(30360) := x"1120";
    tmp(30361) := x"1120";
    tmp(30362) := x"1120";
    tmp(30363) := x"1120";
    tmp(30364) := x"1141";
    tmp(30365) := x"1141";
    tmp(30366) := x"1941";
    tmp(30367) := x"1961";
    tmp(30368) := x"1982";
    tmp(30369) := x"2182";
    tmp(30370) := x"1983";
    tmp(30371) := x"1962";
    tmp(30372) := x"1941";
    tmp(30373) := x"1121";
    tmp(30374) := x"1100";
    tmp(30375) := x"1921";
    tmp(30376) := x"1961";
    tmp(30377) := x"29a1";
    tmp(30378) := x"3a22";
    tmp(30379) := x"4263";
    tmp(30380) := x"4a83";
    tmp(30381) := x"5284";
    tmp(30382) := x"52c5";
    tmp(30383) := x"52a5";
    tmp(30384) := x"5285";
    tmp(30385) := x"5285";
    tmp(30386) := x"5285";
    tmp(30387) := x"5285";
    tmp(30388) := x"4a65";
    tmp(30389) := x"4224";
    tmp(30390) := x"39e3";
    tmp(30391) := x"3182";
    tmp(30392) := x"2122";
    tmp(30393) := x"2121";
    tmp(30394) := x"2121";
    tmp(30395) := x"2141";
    tmp(30396) := x"2962";
    tmp(30397) := x"2962";
    tmp(30398) := x"2982";
    tmp(30399) := x"2982";
    tmp(30400) := x"3182";
    tmp(30401) := x"39c3";
    tmp(30402) := x"4a25";
    tmp(30403) := x"5245";
    tmp(30404) := x"5225";
    tmp(30405) := x"4204";
    tmp(30406) := x"39c4";
    tmp(30407) := x"39a3";
    tmp(30408) := x"3163";
    tmp(30409) := x"2942";
    tmp(30410) := x"2943";
    tmp(30411) := x"2923";
    tmp(30412) := x"2943";
    tmp(30413) := x"3164";
    tmp(30414) := x"3164";
    tmp(30415) := x"3164";
    tmp(30416) := x"3985";
    tmp(30417) := x"39a5";
    tmp(30418) := x"41c6";
    tmp(30419) := x"49c7";
    tmp(30420) := x"49e7";
    tmp(30421) := x"5208";
    tmp(30422) := x"5209";
    tmp(30423) := x"5a4a";
    tmp(30424) := x"6aab";
    tmp(30425) := x"72cd";
    tmp(30426) := x"7b0e";
    tmp(30427) := x"7b2f";
    tmp(30428) := x"8b90";
    tmp(30429) := x"8b91";
    tmp(30430) := x"93d2";
    tmp(30431) := x"93f3";
    tmp(30432) := x"9c14";
    tmp(30433) := x"9c14";
    tmp(30434) := x"9c14";
    tmp(30435) := x"93f4";
    tmp(30436) := x"93d3";
    tmp(30437) := x"07e0";
    tmp(30438) := x"07e0";
    tmp(30439) := x"07e0";
    tmp(30440) := x"07e0";
    tmp(30441) := x"07e0";
    tmp(30442) := x"07e0";
    tmp(30443) := x"07e0";
    tmp(30444) := x"07e0";
    tmp(30445) := x"07e0";
    tmp(30446) := x"07e0";
    tmp(30447) := x"07e0";
    tmp(30448) := x"07e0";
    tmp(30449) := x"07e0";
    tmp(30450) := x"07e0";
    tmp(30451) := x"07e0";
    tmp(30452) := x"07e0";
    tmp(30453) := x"07e0";
    tmp(30454) := x"07e0";
    tmp(30455) := x"07e0";
    tmp(30456) := x"07e0";
    tmp(30457) := x"07e0";
    tmp(30458) := x"07e0";
    tmp(30459) := x"07e0";
    tmp(30460) := x"07e0";
    tmp(30461) := x"07e0";
    tmp(30462) := x"07e0";
    tmp(30463) := x"07e0";
    tmp(30464) := x"07e0";
    tmp(30465) := x"07e0";
    tmp(30466) := x"07e0";
    tmp(30467) := x"07e0";
    tmp(30468) := x"07e0";
    tmp(30469) := x"07e0";
    tmp(30470) := x"07e0";
    tmp(30471) := x"07e0";
    tmp(30472) := x"07e0";
    tmp(30473) := x"07e0";
    tmp(30474) := x"07e0";
    tmp(30475) := x"07e0";
    tmp(30476) := x"07e0";
    tmp(30477) := x"0840";
    tmp(30478) := x"0840";
    tmp(30479) := x"0840";
    tmp(30480) := x"0000";
    tmp(30481) := x"00a4";
    tmp(30482) := x"00a4";
    tmp(30483) := x"00a4";
    tmp(30484) := x"00c4";
    tmp(30485) := x"00c4";
    tmp(30486) := x"00c4";
    tmp(30487) := x"00c5";
    tmp(30488) := x"00c4";
    tmp(30489) := x"00a4";
    tmp(30490) := x"0083";
    tmp(30491) := x"0021";
    tmp(30492) := x"0000";
    tmp(30493) := x"0000";
    tmp(30494) := x"0020";
    tmp(30495) := x"0882";
    tmp(30496) := x"08a3";
    tmp(30497) := x"08a3";
    tmp(30498) := x"08a4";
    tmp(30499) := x"08c4";
    tmp(30500) := x"08c4";
    tmp(30501) := x"08e5";
    tmp(30502) := x"08c5";
    tmp(30503) := x"08c5";
    tmp(30504) := x"08c5";
    tmp(30505) := x"08c5";
    tmp(30506) := x"08c4";
    tmp(30507) := x"08c4";
    tmp(30508) := x"08a4";
    tmp(30509) := x"08a3";
    tmp(30510) := x"0883";
    tmp(30511) := x"0883";
    tmp(30512) := x"08c4";
    tmp(30513) := x"0906";
    tmp(30514) := x"08e5";
    tmp(30515) := x"08c4";
    tmp(30516) := x"08e4";
    tmp(30517) := x"08e5";
    tmp(30518) := x"0926";
    tmp(30519) := x"08e5";
    tmp(30520) := x"08c4";
    tmp(30521) := x"08e5";
    tmp(30522) := x"08e5";
    tmp(30523) := x"0905";
    tmp(30524) := x"0905";
    tmp(30525) := x"0905";
    tmp(30526) := x"08a3";
    tmp(30527) := x"0062";
    tmp(30528) := x"0882";
    tmp(30529) := x"08c4";
    tmp(30530) := x"0905";
    tmp(30531) := x"0905";
    tmp(30532) := x"0905";
    tmp(30533) := x"0905";
    tmp(30534) := x"0904";
    tmp(30535) := x"0905";
    tmp(30536) := x"1104";
    tmp(30537) := x"08a3";
    tmp(30538) := x"0861";
    tmp(30539) := x"10e3";
    tmp(30540) := x"1124";
    tmp(30541) := x"08c1";
    tmp(30542) := x"08c0";
    tmp(30543) := x"08c0";
    tmp(30544) := x"08c0";
    tmp(30545) := x"08c0";
    tmp(30546) := x"08c0";
    tmp(30547) := x"08c0";
    tmp(30548) := x"08c0";
    tmp(30549) := x"08e0";
    tmp(30550) := x"1101";
    tmp(30551) := x"1121";
    tmp(30552) := x"1962";
    tmp(30553) := x"21a3";
    tmp(30554) := x"31e4";
    tmp(30555) := x"3a25";
    tmp(30556) := x"4a87";
    tmp(30557) := x"52a9";
    tmp(30558) := x"6b2b";
    tmp(30559) := x"7bad";
    tmp(30560) := x"8c10";
    tmp(30561) := x"9451";
    tmp(30562) := x"9472";
    tmp(30563) := x"9493";
    tmp(30564) := x"9494";
    tmp(30565) := x"9cb6";
    tmp(30566) := x"a4d7";
    tmp(30567) := x"a4d7";
    tmp(30568) := x"9497";
    tmp(30569) := x"a518";
    tmp(30570) := x"9cd8";
    tmp(30571) := x"9cd8";
    tmp(30572) := x"9cf9";
    tmp(30573) := x"9d19";
    tmp(30574) := x"94f9";
    tmp(30575) := x"94d9";
    tmp(30576) := x"94d9";
    tmp(30577) := x"8cb7";
    tmp(30578) := x"8455";
    tmp(30579) := x"8453";
    tmp(30580) := x"7c11";
    tmp(30581) := x"73ce";
    tmp(30582) := x"6b8c";
    tmp(30583) := x"5b0a";
    tmp(30584) := x"52c7";
    tmp(30585) := x"4265";
    tmp(30586) := x"3204";
    tmp(30587) := x"21c3";
    tmp(30588) := x"1982";
    tmp(30589) := x"1162";
    tmp(30590) := x"1162";
    tmp(30591) := x"1183";
    tmp(30592) := x"1183";
    tmp(30593) := x"19c3";
    tmp(30594) := x"2203";
    tmp(30595) := x"2a24";
    tmp(30596) := x"3263";
    tmp(30597) := x"2202";
    tmp(30598) := x"1141";
    tmp(30599) := x"1121";
    tmp(30600) := x"1121";
    tmp(30601) := x"1121";
    tmp(30602) := x"1120";
    tmp(30603) := x"1120";
    tmp(30604) := x"1120";
    tmp(30605) := x"1141";
    tmp(30606) := x"1941";
    tmp(30607) := x"1941";
    tmp(30608) := x"1962";
    tmp(30609) := x"2183";
    tmp(30610) := x"21a3";
    tmp(30611) := x"1962";
    tmp(30612) := x"1941";
    tmp(30613) := x"1121";
    tmp(30614) := x"1100";
    tmp(30615) := x"1120";
    tmp(30616) := x"1941";
    tmp(30617) := x"2161";
    tmp(30618) := x"29c1";
    tmp(30619) := x"3202";
    tmp(30620) := x"4243";
    tmp(30621) := x"4264";
    tmp(30622) := x"4a64";
    tmp(30623) := x"4a84";
    tmp(30624) := x"4a84";
    tmp(30625) := x"4a85";
    tmp(30626) := x"4a44";
    tmp(30627) := x"4a65";
    tmp(30628) := x"4224";
    tmp(30629) := x"4224";
    tmp(30630) := x"4204";
    tmp(30631) := x"31a3";
    tmp(30632) := x"2962";
    tmp(30633) := x"2121";
    tmp(30634) := x"2121";
    tmp(30635) := x"2141";
    tmp(30636) := x"2962";
    tmp(30637) := x"2982";
    tmp(30638) := x"2982";
    tmp(30639) := x"2982";
    tmp(30640) := x"2962";
    tmp(30641) := x"3183";
    tmp(30642) := x"39c3";
    tmp(30643) := x"41e4";
    tmp(30644) := x"4a04";
    tmp(30645) := x"41c4";
    tmp(30646) := x"39a3";
    tmp(30647) := x"3183";
    tmp(30648) := x"2942";
    tmp(30649) := x"2922";
    tmp(30650) := x"2922";
    tmp(30651) := x"2923";
    tmp(30652) := x"2943";
    tmp(30653) := x"3143";
    tmp(30654) := x"3164";
    tmp(30655) := x"3164";
    tmp(30656) := x"3164";
    tmp(30657) := x"39a5";
    tmp(30658) := x"39a5";
    tmp(30659) := x"41a6";
    tmp(30660) := x"41a6";
    tmp(30661) := x"49c7";
    tmp(30662) := x"5208";
    tmp(30663) := x"5228";
    tmp(30664) := x"624a";
    tmp(30665) := x"6a8b";
    tmp(30666) := x"6aad";
    tmp(30667) := x"72ee";
    tmp(30668) := x"7b0f";
    tmp(30669) := x"834f";
    tmp(30670) := x"8371";
    tmp(30671) := x"8b91";
    tmp(30672) := x"8bb2";
    tmp(30673) := x"93f3";
    tmp(30674) := x"8bb2";
    tmp(30675) := x"8bb2";
    tmp(30676) := x"93d2";
    tmp(30677) := x"07e0";
    tmp(30678) := x"07e0";
    tmp(30679) := x"07e0";
    tmp(30680) := x"07e0";
    tmp(30681) := x"07e0";
    tmp(30682) := x"07e0";
    tmp(30683) := x"07e0";
    tmp(30684) := x"07e0";
    tmp(30685) := x"07e0";
    tmp(30686) := x"07e0";
    tmp(30687) := x"07e0";
    tmp(30688) := x"07e0";
    tmp(30689) := x"07e0";
    tmp(30690) := x"07e0";
    tmp(30691) := x"07e0";
    tmp(30692) := x"07e0";
    tmp(30693) := x"07e0";
    tmp(30694) := x"07e0";
    tmp(30695) := x"07e0";
    tmp(30696) := x"07e0";
    tmp(30697) := x"07e0";
    tmp(30698) := x"07e0";
    tmp(30699) := x"07e0";
    tmp(30700) := x"07e0";
    tmp(30701) := x"07e0";
    tmp(30702) := x"07e0";
    tmp(30703) := x"07e0";
    tmp(30704) := x"07e0";
    tmp(30705) := x"07e0";
    tmp(30706) := x"07e0";
    tmp(30707) := x"07e0";
    tmp(30708) := x"07e0";
    tmp(30709) := x"07e0";
    tmp(30710) := x"07e0";
    tmp(30711) := x"07e0";
    tmp(30712) := x"07e0";
    tmp(30713) := x"07e0";
    tmp(30714) := x"07e0";
    tmp(30715) := x"07e0";
    tmp(30716) := x"07e0";
    tmp(30717) := x"0840";
    tmp(30718) := x"0840";
    tmp(30719) := x"0840";
    tmp(30720) := x"0000";
    tmp(30721) := x"00a4";
    tmp(30722) := x"00a4";
    tmp(30723) := x"00c4";
    tmp(30724) := x"00a4";
    tmp(30725) := x"00c4";
    tmp(30726) := x"00c4";
    tmp(30727) := x"00c4";
    tmp(30728) := x"00c4";
    tmp(30729) := x"0062";
    tmp(30730) := x"0041";
    tmp(30731) := x"0021";
    tmp(30732) := x"0020";
    tmp(30733) := x"0000";
    tmp(30734) := x"0021";
    tmp(30735) := x"0862";
    tmp(30736) := x"0882";
    tmp(30737) := x"08a3";
    tmp(30738) := x"08a4";
    tmp(30739) := x"0883";
    tmp(30740) := x"0062";
    tmp(30741) := x"08a3";
    tmp(30742) := x"08c4";
    tmp(30743) := x"08a4";
    tmp(30744) := x"08a4";
    tmp(30745) := x"08a4";
    tmp(30746) := x"08a4";
    tmp(30747) := x"08a4";
    tmp(30748) := x"08a4";
    tmp(30749) := x"08a4";
    tmp(30750) := x"08c5";
    tmp(30751) := x"0905";
    tmp(30752) := x"0905";
    tmp(30753) := x"08e5";
    tmp(30754) := x"0926";
    tmp(30755) := x"0905";
    tmp(30756) := x"0905";
    tmp(30757) := x"0905";
    tmp(30758) := x"08e5";
    tmp(30759) := x"0905";
    tmp(30760) := x"08e5";
    tmp(30761) := x"08e4";
    tmp(30762) := x"08c4";
    tmp(30763) := x"08e5";
    tmp(30764) := x"0905";
    tmp(30765) := x"08e4";
    tmp(30766) := x"0882";
    tmp(30767) := x"0062";
    tmp(30768) := x"08c3";
    tmp(30769) := x"0905";
    tmp(30770) := x"08e4";
    tmp(30771) := x"0904";
    tmp(30772) := x"08e4";
    tmp(30773) := x"08c4";
    tmp(30774) := x"08c4";
    tmp(30775) := x"08c3";
    tmp(30776) := x"08c3";
    tmp(30777) := x"08c3";
    tmp(30778) := x"08e3";
    tmp(30779) := x"1104";
    tmp(30780) := x"08a1";
    tmp(30781) := x"08c1";
    tmp(30782) := x"08e0";
    tmp(30783) := x"08e0";
    tmp(30784) := x"08e0";
    tmp(30785) := x"08e0";
    tmp(30786) := x"08e0";
    tmp(30787) := x"08e0";
    tmp(30788) := x"08e0";
    tmp(30789) := x"08e0";
    tmp(30790) := x"08e0";
    tmp(30791) := x"1101";
    tmp(30792) := x"1941";
    tmp(30793) := x"2182";
    tmp(30794) := x"29a3";
    tmp(30795) := x"3204";
    tmp(30796) := x"4246";
    tmp(30797) := x"4a88";
    tmp(30798) := x"5aea";
    tmp(30799) := x"632b";
    tmp(30800) := x"736d";
    tmp(30801) := x"7bae";
    tmp(30802) := x"8411";
    tmp(30803) := x"8c31";
    tmp(30804) := x"8c32";
    tmp(30805) := x"9453";
    tmp(30806) := x"9454";
    tmp(30807) := x"9c76";
    tmp(30808) := x"9456";
    tmp(30809) := x"9496";
    tmp(30810) := x"9476";
    tmp(30811) := x"9497";
    tmp(30812) := x"8c56";
    tmp(30813) := x"94b7";
    tmp(30814) := x"8c97";
    tmp(30815) := x"8c76";
    tmp(30816) := x"8455";
    tmp(30817) := x"7c34";
    tmp(30818) := x"73f2";
    tmp(30819) := x"73d0";
    tmp(30820) := x"6b8e";
    tmp(30821) := x"636c";
    tmp(30822) := x"5b09";
    tmp(30823) := x"4aa7";
    tmp(30824) := x"4245";
    tmp(30825) := x"3204";
    tmp(30826) := x"29a3";
    tmp(30827) := x"2183";
    tmp(30828) := x"1962";
    tmp(30829) := x"1163";
    tmp(30830) := x"1163";
    tmp(30831) := x"1183";
    tmp(30832) := x"19a3";
    tmp(30833) := x"21c3";
    tmp(30834) := x"2a03";
    tmp(30835) := x"3244";
    tmp(30836) := x"2a43";
    tmp(30837) := x"19a1";
    tmp(30838) := x"1121";
    tmp(30839) := x"1121";
    tmp(30840) := x"1121";
    tmp(30841) := x"1121";
    tmp(30842) := x"1121";
    tmp(30843) := x"1120";
    tmp(30844) := x"1120";
    tmp(30845) := x"1120";
    tmp(30846) := x"1141";
    tmp(30847) := x"1941";
    tmp(30848) := x"1962";
    tmp(30849) := x"2182";
    tmp(30850) := x"21a3";
    tmp(30851) := x"1982";
    tmp(30852) := x"1941";
    tmp(30853) := x"1121";
    tmp(30854) := x"1101";
    tmp(30855) := x"1120";
    tmp(30856) := x"1940";
    tmp(30857) := x"1961";
    tmp(30858) := x"2181";
    tmp(30859) := x"29c1";
    tmp(30860) := x"3202";
    tmp(30861) := x"4223";
    tmp(30862) := x"4243";
    tmp(30863) := x"4a44";
    tmp(30864) := x"4244";
    tmp(30865) := x"4a44";
    tmp(30866) := x"4224";
    tmp(30867) := x"4224";
    tmp(30868) := x"4224";
    tmp(30869) := x"4224";
    tmp(30870) := x"39e3";
    tmp(30871) := x"39e3";
    tmp(30872) := x"3183";
    tmp(30873) := x"2942";
    tmp(30874) := x"2122";
    tmp(30875) := x"2142";
    tmp(30876) := x"2142";
    tmp(30877) := x"2962";
    tmp(30878) := x"2962";
    tmp(30879) := x"2982";
    tmp(30880) := x"2962";
    tmp(30881) := x"2982";
    tmp(30882) := x"3183";
    tmp(30883) := x"39a3";
    tmp(30884) := x"41c4";
    tmp(30885) := x"39c4";
    tmp(30886) := x"3183";
    tmp(30887) := x"2962";
    tmp(30888) := x"2942";
    tmp(30889) := x"2922";
    tmp(30890) := x"2922";
    tmp(30891) := x"2923";
    tmp(30892) := x"2923";
    tmp(30893) := x"2943";
    tmp(30894) := x"3143";
    tmp(30895) := x"3144";
    tmp(30896) := x"3164";
    tmp(30897) := x"3144";
    tmp(30898) := x"3965";
    tmp(30899) := x"4185";
    tmp(30900) := x"41a6";
    tmp(30901) := x"41a6";
    tmp(30902) := x"49e7";
    tmp(30903) := x"51e8";
    tmp(30904) := x"5a08";
    tmp(30905) := x"624a";
    tmp(30906) := x"626b";
    tmp(30907) := x"6a8b";
    tmp(30908) := x"6aac";
    tmp(30909) := x"72ed";
    tmp(30910) := x"730e";
    tmp(30911) := x"7b0e";
    tmp(30912) := x"834f";
    tmp(30913) := x"8350";
    tmp(30914) := x"8350";
    tmp(30915) := x"8371";
    tmp(30916) := x"7b50";
    tmp(30917) := x"07e0";
    tmp(30918) := x"07e0";
    tmp(30919) := x"07e0";
    tmp(30920) := x"07e0";
    tmp(30921) := x"07e0";
    tmp(30922) := x"07e0";
    tmp(30923) := x"07e0";
    tmp(30924) := x"07e0";
    tmp(30925) := x"07e0";
    tmp(30926) := x"07e0";
    tmp(30927) := x"07e0";
    tmp(30928) := x"07e0";
    tmp(30929) := x"07e0";
    tmp(30930) := x"07e0";
    tmp(30931) := x"07e0";
    tmp(30932) := x"07e0";
    tmp(30933) := x"07e0";
    tmp(30934) := x"07e0";
    tmp(30935) := x"07e0";
    tmp(30936) := x"07e0";
    tmp(30937) := x"07e0";
    tmp(30938) := x"07e0";
    tmp(30939) := x"07e0";
    tmp(30940) := x"07e0";
    tmp(30941) := x"07e0";
    tmp(30942) := x"07e0";
    tmp(30943) := x"07e0";
    tmp(30944) := x"07e0";
    tmp(30945) := x"07e0";
    tmp(30946) := x"07e0";
    tmp(30947) := x"07e0";
    tmp(30948) := x"07e0";
    tmp(30949) := x"07e0";
    tmp(30950) := x"07e0";
    tmp(30951) := x"07e0";
    tmp(30952) := x"07e0";
    tmp(30953) := x"07e0";
    tmp(30954) := x"07e0";
    tmp(30955) := x"07e0";
    tmp(30956) := x"07e0";
    tmp(30957) := x"0840";
    tmp(30958) := x"0840";
    tmp(30959) := x"0840";
    tmp(30960) := x"0020";
    tmp(30961) := x"00c4";
    tmp(30962) := x"00c4";
    tmp(30963) := x"00c4";
    tmp(30964) := x"00a4";
    tmp(30965) := x"00c4";
    tmp(30966) := x"00a4";
    tmp(30967) := x"00a4";
    tmp(30968) := x"00a4";
    tmp(30969) := x"0041";
    tmp(30970) := x"0041";
    tmp(30971) := x"0021";
    tmp(30972) := x"0020";
    tmp(30973) := x"0021";
    tmp(30974) := x"0841";
    tmp(30975) := x"0862";
    tmp(30976) := x"08a3";
    tmp(30977) := x"0882";
    tmp(30978) := x"08a3";
    tmp(30979) := x"0883";
    tmp(30980) := x"08a3";
    tmp(30981) := x"08a3";
    tmp(30982) := x"08a3";
    tmp(30983) := x"08a3";
    tmp(30984) := x"08a3";
    tmp(30985) := x"0883";
    tmp(30986) := x"08a3";
    tmp(30987) := x"0083";
    tmp(30988) := x"08a4";
    tmp(30989) := x"08e5";
    tmp(30990) := x"0905";
    tmp(30991) := x"08e5";
    tmp(30992) := x"08e4";
    tmp(30993) := x"08c4";
    tmp(30994) := x"00c4";
    tmp(30995) := x"0905";
    tmp(30996) := x"0925";
    tmp(30997) := x"08e4";
    tmp(30998) := x"08c4";
    tmp(30999) := x"0905";
    tmp(31000) := x"08e5";
    tmp(31001) := x"0905";
    tmp(31002) := x"0946";
    tmp(31003) := x"0926";
    tmp(31004) := x"0905";
    tmp(31005) := x"0925";
    tmp(31006) := x"08e4";
    tmp(31007) := x"0904";
    tmp(31008) := x"0925";
    tmp(31009) := x"0925";
    tmp(31010) := x"0905";
    tmp(31011) := x"08e4";
    tmp(31012) := x"08e4";
    tmp(31013) := x"08e4";
    tmp(31014) := x"1125";
    tmp(31015) := x"1105";
    tmp(31016) := x"1125";
    tmp(31017) := x"1104";
    tmp(31018) := x"08c3";
    tmp(31019) := x"0881";
    tmp(31020) := x"10e1";
    tmp(31021) := x"08e0";
    tmp(31022) := x"0900";
    tmp(31023) := x"0900";
    tmp(31024) := x"08e0";
    tmp(31025) := x"08e0";
    tmp(31026) := x"08e0";
    tmp(31027) := x"08e0";
    tmp(31028) := x"08e0";
    tmp(31029) := x"08e0";
    tmp(31030) := x"0900";
    tmp(31031) := x"0901";
    tmp(31032) := x"1121";
    tmp(31033) := x"1942";
    tmp(31034) := x"2182";
    tmp(31035) := x"29c4";
    tmp(31036) := x"3205";
    tmp(31037) := x"3a46";
    tmp(31038) := x"4a88";
    tmp(31039) := x"5aca";
    tmp(31040) := x"6b4b";
    tmp(31041) := x"6b6d";
    tmp(31042) := x"736d";
    tmp(31043) := x"83af";
    tmp(31044) := x"7bb0";
    tmp(31045) := x"7bb1";
    tmp(31046) := x"83d2";
    tmp(31047) := x"83f2";
    tmp(31048) := x"8413";
    tmp(31049) := x"7bf3";
    tmp(31050) := x"8434";
    tmp(31051) := x"83d3";
    tmp(31052) := x"8c55";
    tmp(31053) := x"8c75";
    tmp(31054) := x"8434";
    tmp(31055) := x"8414";
    tmp(31056) := x"73f2";
    tmp(31057) := x"73f1";
    tmp(31058) := x"6b8e";
    tmp(31059) := x"636d";
    tmp(31060) := x"634b";
    tmp(31061) := x"52e9";
    tmp(31062) := x"4ac7";
    tmp(31063) := x"4266";
    tmp(31064) := x"3204";
    tmp(31065) := x"29a3";
    tmp(31066) := x"21a3";
    tmp(31067) := x"1963";
    tmp(31068) := x"1963";
    tmp(31069) := x"1163";
    tmp(31070) := x"1163";
    tmp(31071) := x"1983";
    tmp(31072) := x"19a3";
    tmp(31073) := x"21e4";
    tmp(31074) := x"2a24";
    tmp(31075) := x"2a43";
    tmp(31076) := x"2202";
    tmp(31077) := x"1161";
    tmp(31078) := x"1121";
    tmp(31079) := x"1121";
    tmp(31080) := x"1141";
    tmp(31081) := x"1121";
    tmp(31082) := x"1121";
    tmp(31083) := x"1120";
    tmp(31084) := x"1120";
    tmp(31085) := x"1120";
    tmp(31086) := x"1141";
    tmp(31087) := x"1941";
    tmp(31088) := x"1961";
    tmp(31089) := x"2182";
    tmp(31090) := x"21a2";
    tmp(31091) := x"1982";
    tmp(31092) := x"1941";
    tmp(31093) := x"1121";
    tmp(31094) := x"1121";
    tmp(31095) := x"1100";
    tmp(31096) := x"1920";
    tmp(31097) := x"1941";
    tmp(31098) := x"1941";
    tmp(31099) := x"2181";
    tmp(31100) := x"29c1";
    tmp(31101) := x"3202";
    tmp(31102) := x"3a23";
    tmp(31103) := x"3a23";
    tmp(31104) := x"4223";
    tmp(31105) := x"4224";
    tmp(31106) := x"4204";
    tmp(31107) := x"4204";
    tmp(31108) := x"4224";
    tmp(31109) := x"39e4";
    tmp(31110) := x"39e3";
    tmp(31111) := x"39c3";
    tmp(31112) := x"31a3";
    tmp(31113) := x"2962";
    tmp(31114) := x"2942";
    tmp(31115) := x"2942";
    tmp(31116) := x"2962";
    tmp(31117) := x"2962";
    tmp(31118) := x"2962";
    tmp(31119) := x"2982";
    tmp(31120) := x"2982";
    tmp(31121) := x"2982";
    tmp(31122) := x"2983";
    tmp(31123) := x"3183";
    tmp(31124) := x"31a3";
    tmp(31125) := x"31a3";
    tmp(31126) := x"3183";
    tmp(31127) := x"2962";
    tmp(31128) := x"2942";
    tmp(31129) := x"2922";
    tmp(31130) := x"2922";
    tmp(31131) := x"2922";
    tmp(31132) := x"2923";
    tmp(31133) := x"2943";
    tmp(31134) := x"2923";
    tmp(31135) := x"2923";
    tmp(31136) := x"3144";
    tmp(31137) := x"3164";
    tmp(31138) := x"3144";
    tmp(31139) := x"3965";
    tmp(31140) := x"3985";
    tmp(31141) := x"41a6";
    tmp(31142) := x"41a6";
    tmp(31143) := x"49a7";
    tmp(31144) := x"51e7";
    tmp(31145) := x"51e8";
    tmp(31146) := x"5208";
    tmp(31147) := x"5a49";
    tmp(31148) := x"626a";
    tmp(31149) := x"628b";
    tmp(31150) := x"6aac";
    tmp(31151) := x"6acc";
    tmp(31152) := x"72ed";
    tmp(31153) := x"72ed";
    tmp(31154) := x"6aed";
    tmp(31155) := x"730e";
    tmp(31156) := x"730e";
    tmp(31157) := x"07e0";
    tmp(31158) := x"07e0";
    tmp(31159) := x"07e0";
    tmp(31160) := x"07e0";
    tmp(31161) := x"07e0";
    tmp(31162) := x"07e0";
    tmp(31163) := x"07e0";
    tmp(31164) := x"07e0";
    tmp(31165) := x"07e0";
    tmp(31166) := x"07e0";
    tmp(31167) := x"07e0";
    tmp(31168) := x"07e0";
    tmp(31169) := x"07e0";
    tmp(31170) := x"07e0";
    tmp(31171) := x"07e0";
    tmp(31172) := x"07e0";
    tmp(31173) := x"07e0";
    tmp(31174) := x"07e0";
    tmp(31175) := x"07e0";
    tmp(31176) := x"07e0";
    tmp(31177) := x"07e0";
    tmp(31178) := x"07e0";
    tmp(31179) := x"07e0";
    tmp(31180) := x"07e0";
    tmp(31181) := x"07e0";
    tmp(31182) := x"07e0";
    tmp(31183) := x"07e0";
    tmp(31184) := x"07e0";
    tmp(31185) := x"07e0";
    tmp(31186) := x"07e0";
    tmp(31187) := x"07e0";
    tmp(31188) := x"07e0";
    tmp(31189) := x"07e0";
    tmp(31190) := x"07e0";
    tmp(31191) := x"07e0";
    tmp(31192) := x"07e0";
    tmp(31193) := x"07e0";
    tmp(31194) := x"07e0";
    tmp(31195) := x"07e0";
    tmp(31196) := x"07e0";
    tmp(31197) := x"0840";
    tmp(31198) := x"0840";
    tmp(31199) := x"0840";
    tmp(31200) := x"0020";
    tmp(31201) := x"00c4";
    tmp(31202) := x"00c4";
    tmp(31203) := x"00a4";
    tmp(31204) := x"00a4";
    tmp(31205) := x"00a4";
    tmp(31206) := x"00a4";
    tmp(31207) := x"00a4";
    tmp(31208) := x"00a3";
    tmp(31209) := x"0062";
    tmp(31210) := x"0062";
    tmp(31211) := x"0082";
    tmp(31212) := x"0021";
    tmp(31213) := x"0021";
    tmp(31214) := x"0041";
    tmp(31215) := x"0062";
    tmp(31216) := x"0882";
    tmp(31217) := x"0882";
    tmp(31218) := x"0882";
    tmp(31219) := x"0882";
    tmp(31220) := x"08a3";
    tmp(31221) := x"08a3";
    tmp(31222) := x"08a3";
    tmp(31223) := x"08a3";
    tmp(31224) := x"0883";
    tmp(31225) := x"0883";
    tmp(31226) := x"00a3";
    tmp(31227) := x"0905";
    tmp(31228) := x"0906";
    tmp(31229) := x"0905";
    tmp(31230) := x"08e5";
    tmp(31231) := x"08e4";
    tmp(31232) := x"08e4";
    tmp(31233) := x"08c4";
    tmp(31234) := x"0905";
    tmp(31235) := x"0926";
    tmp(31236) := x"0905";
    tmp(31237) := x"08e5";
    tmp(31238) := x"0905";
    tmp(31239) := x"0905";
    tmp(31240) := x"0906";
    tmp(31241) := x"0947";
    tmp(31242) := x"0947";
    tmp(31243) := x"0926";
    tmp(31244) := x"0926";
    tmp(31245) := x"0926";
    tmp(31246) := x"0925";
    tmp(31247) := x"0925";
    tmp(31248) := x"08e4";
    tmp(31249) := x"08c3";
    tmp(31250) := x"08c3";
    tmp(31251) := x"0904";
    tmp(31252) := x"08c3";
    tmp(31253) := x"08c3";
    tmp(31254) := x"08e3";
    tmp(31255) := x"08c3";
    tmp(31256) := x"08a3";
    tmp(31257) := x"08a3";
    tmp(31258) := x"0861";
    tmp(31259) := x"08a1";
    tmp(31260) := x"0901";
    tmp(31261) := x"0900";
    tmp(31262) := x"0900";
    tmp(31263) := x"0900";
    tmp(31264) := x"0900";
    tmp(31265) := x"0900";
    tmp(31266) := x"0900";
    tmp(31267) := x"0900";
    tmp(31268) := x"0900";
    tmp(31269) := x"08e0";
    tmp(31270) := x"08e0";
    tmp(31271) := x"0900";
    tmp(31272) := x"1101";
    tmp(31273) := x"1121";
    tmp(31274) := x"1962";
    tmp(31275) := x"21a3";
    tmp(31276) := x"31e4";
    tmp(31277) := x"3a25";
    tmp(31278) := x"4247";
    tmp(31279) := x"4a89";
    tmp(31280) := x"5aca";
    tmp(31281) := x"5aeb";
    tmp(31282) := x"632c";
    tmp(31283) := x"6b4e";
    tmp(31284) := x"736e";
    tmp(31285) := x"736f";
    tmp(31286) := x"6b4f";
    tmp(31287) := x"7bb1";
    tmp(31288) := x"7bb1";
    tmp(31289) := x"7bb1";
    tmp(31290) := x"7bb2";
    tmp(31291) := x"7bf3";
    tmp(31292) := x"7bd3";
    tmp(31293) := x"73b2";
    tmp(31294) := x"7bd2";
    tmp(31295) := x"7391";
    tmp(31296) := x"6b6f";
    tmp(31297) := x"634d";
    tmp(31298) := x"632c";
    tmp(31299) := x"5b0b";
    tmp(31300) := x"52c9";
    tmp(31301) := x"4a87";
    tmp(31302) := x"4246";
    tmp(31303) := x"3a04";
    tmp(31304) := x"29a3";
    tmp(31305) := x"2183";
    tmp(31306) := x"2163";
    tmp(31307) := x"1963";
    tmp(31308) := x"1983";
    tmp(31309) := x"1963";
    tmp(31310) := x"1983";
    tmp(31311) := x"19a3";
    tmp(31312) := x"21c3";
    tmp(31313) := x"2a04";
    tmp(31314) := x"2a23";
    tmp(31315) := x"2a22";
    tmp(31316) := x"19a1";
    tmp(31317) := x"1141";
    tmp(31318) := x"1121";
    tmp(31319) := x"1121";
    tmp(31320) := x"1121";
    tmp(31321) := x"1121";
    tmp(31322) := x"1121";
    tmp(31323) := x"1120";
    tmp(31324) := x"1120";
    tmp(31325) := x"1120";
    tmp(31326) := x"1120";
    tmp(31327) := x"1941";
    tmp(31328) := x"1961";
    tmp(31329) := x"1962";
    tmp(31330) := x"2182";
    tmp(31331) := x"1982";
    tmp(31332) := x"1941";
    tmp(31333) := x"1121";
    tmp(31334) := x"1101";
    tmp(31335) := x"1120";
    tmp(31336) := x"1920";
    tmp(31337) := x"1941";
    tmp(31338) := x"1941";
    tmp(31339) := x"2161";
    tmp(31340) := x"2181";
    tmp(31341) := x"29c1";
    tmp(31342) := x"31e2";
    tmp(31343) := x"3a02";
    tmp(31344) := x"3a03";
    tmp(31345) := x"3a23";
    tmp(31346) := x"3a03";
    tmp(31347) := x"39e3";
    tmp(31348) := x"3a03";
    tmp(31349) := x"39e3";
    tmp(31350) := x"31a3";
    tmp(31351) := x"31a3";
    tmp(31352) := x"3183";
    tmp(31353) := x"31a2";
    tmp(31354) := x"2942";
    tmp(31355) := x"2942";
    tmp(31356) := x"2942";
    tmp(31357) := x"2942";
    tmp(31358) := x"2962";
    tmp(31359) := x"2982";
    tmp(31360) := x"2962";
    tmp(31361) := x"2962";
    tmp(31362) := x"2962";
    tmp(31363) := x"2963";
    tmp(31364) := x"3163";
    tmp(31365) := x"3183";
    tmp(31366) := x"3163";
    tmp(31367) := x"2942";
    tmp(31368) := x"2942";
    tmp(31369) := x"2942";
    tmp(31370) := x"2122";
    tmp(31371) := x"2902";
    tmp(31372) := x"2923";
    tmp(31373) := x"2923";
    tmp(31374) := x"2923";
    tmp(31375) := x"2923";
    tmp(31376) := x"2923";
    tmp(31377) := x"3123";
    tmp(31378) := x"3144";
    tmp(31379) := x"3965";
    tmp(31380) := x"3965";
    tmp(31381) := x"3965";
    tmp(31382) := x"3965";
    tmp(31383) := x"4186";
    tmp(31384) := x"41a6";
    tmp(31385) := x"49c6";
    tmp(31386) := x"49c7";
    tmp(31387) := x"49c7";
    tmp(31388) := x"51e8";
    tmp(31389) := x"5229";
    tmp(31390) := x"5a29";
    tmp(31391) := x"5a4a";
    tmp(31392) := x"626a";
    tmp(31393) := x"626a";
    tmp(31394) := x"628b";
    tmp(31395) := x"628b";
    tmp(31396) := x"5a6b";
    tmp(31397) := x"07e0";
    tmp(31398) := x"07e0";
    tmp(31399) := x"07e0";
    tmp(31400) := x"07e0";
    tmp(31401) := x"07e0";
    tmp(31402) := x"07e0";
    tmp(31403) := x"07e0";
    tmp(31404) := x"07e0";
    tmp(31405) := x"07e0";
    tmp(31406) := x"07e0";
    tmp(31407) := x"07e0";
    tmp(31408) := x"07e0";
    tmp(31409) := x"07e0";
    tmp(31410) := x"07e0";
    tmp(31411) := x"07e0";
    tmp(31412) := x"07e0";
    tmp(31413) := x"07e0";
    tmp(31414) := x"07e0";
    tmp(31415) := x"07e0";
    tmp(31416) := x"07e0";
    tmp(31417) := x"07e0";
    tmp(31418) := x"07e0";
    tmp(31419) := x"07e0";
    tmp(31420) := x"07e0";
    tmp(31421) := x"07e0";
    tmp(31422) := x"07e0";
    tmp(31423) := x"07e0";
    tmp(31424) := x"07e0";
    tmp(31425) := x"07e0";
    tmp(31426) := x"07e0";
    tmp(31427) := x"07e0";
    tmp(31428) := x"07e0";
    tmp(31429) := x"07e0";
    tmp(31430) := x"07e0";
    tmp(31431) := x"07e0";
    tmp(31432) := x"07e0";
    tmp(31433) := x"07e0";
    tmp(31434) := x"07e0";
    tmp(31435) := x"07e0";
    tmp(31436) := x"07e0";
    tmp(31437) := x"0840";
    tmp(31438) := x"0840";
    tmp(31439) := x"0840";
    tmp(31440) := x"0020";
    tmp(31441) := x"00e5";
    tmp(31442) := x"00e5";
    tmp(31443) := x"00c5";
    tmp(31444) := x"00c4";
    tmp(31445) := x"00a4";
    tmp(31446) := x"00a4";
    tmp(31447) := x"00a4";
    tmp(31448) := x"00a4";
    tmp(31449) := x"00a3";
    tmp(31450) := x"0083";
    tmp(31451) := x"0083";
    tmp(31452) := x"0062";
    tmp(31453) := x"0021";
    tmp(31454) := x"0021";
    tmp(31455) := x"0041";
    tmp(31456) := x"0862";
    tmp(31457) := x"0062";
    tmp(31458) := x"08a3";
    tmp(31459) := x"08a3";
    tmp(31460) := x"08a3";
    tmp(31461) := x"0883";
    tmp(31462) := x"0882";
    tmp(31463) := x"0882";
    tmp(31464) := x"0082";
    tmp(31465) := x"08a4";
    tmp(31466) := x"0926";
    tmp(31467) := x"0926";
    tmp(31468) := x"0905";
    tmp(31469) := x"08e5";
    tmp(31470) := x"08e4";
    tmp(31471) := x"08e4";
    tmp(31472) := x"08e4";
    tmp(31473) := x"0905";
    tmp(31474) := x"0926";
    tmp(31475) := x"0905";
    tmp(31476) := x"0905";
    tmp(31477) := x"0905";
    tmp(31478) := x"08e5";
    tmp(31479) := x"08c4";
    tmp(31480) := x"08c5";
    tmp(31481) := x"0906";
    tmp(31482) := x"0926";
    tmp(31483) := x"0925";
    tmp(31484) := x"0905";
    tmp(31485) := x"0904";
    tmp(31486) := x"08e4";
    tmp(31487) := x"08e4";
    tmp(31488) := x"08c3";
    tmp(31489) := x"08c3";
    tmp(31490) := x"0904";
    tmp(31491) := x"0904";
    tmp(31492) := x"08e3";
    tmp(31493) := x"08c3";
    tmp(31494) := x"08c3";
    tmp(31495) := x"08a3";
    tmp(31496) := x"08e3";
    tmp(31497) := x"10c3";
    tmp(31498) := x"08c2";
    tmp(31499) := x"1121";
    tmp(31500) := x"1100";
    tmp(31501) := x"0900";
    tmp(31502) := x"0920";
    tmp(31503) := x"0900";
    tmp(31504) := x"0920";
    tmp(31505) := x"0900";
    tmp(31506) := x"0900";
    tmp(31507) := x"0900";
    tmp(31508) := x"0900";
    tmp(31509) := x"0900";
    tmp(31510) := x"08e0";
    tmp(31511) := x"0900";
    tmp(31512) := x"0901";
    tmp(31513) := x"1121";
    tmp(31514) := x"1941";
    tmp(31515) := x"2182";
    tmp(31516) := x"21a3";
    tmp(31517) := x"29c4";
    tmp(31518) := x"3205";
    tmp(31519) := x"3a47";
    tmp(31520) := x"4a68";
    tmp(31521) := x"52a9";
    tmp(31522) := x"5aeb";
    tmp(31523) := x"630c";
    tmp(31524) := x"630c";
    tmp(31525) := x"6b2d";
    tmp(31526) := x"6b2e";
    tmp(31527) := x"6b2e";
    tmp(31528) := x"6b0e";
    tmp(31529) := x"7350";
    tmp(31530) := x"7351";
    tmp(31531) := x"7371";
    tmp(31532) := x"7372";
    tmp(31533) := x"6b51";
    tmp(31534) := x"6b50";
    tmp(31535) := x"6b2e";
    tmp(31536) := x"630d";
    tmp(31537) := x"630c";
    tmp(31538) := x"5aea";
    tmp(31539) := x"52c9";
    tmp(31540) := x"4a67";
    tmp(31541) := x"4246";
    tmp(31542) := x"3a05";
    tmp(31543) := x"29c4";
    tmp(31544) := x"2983";
    tmp(31545) := x"2183";
    tmp(31546) := x"2163";
    tmp(31547) := x"1984";
    tmp(31548) := x"19a4";
    tmp(31549) := x"1963";
    tmp(31550) := x"1983";
    tmp(31551) := x"19a3";
    tmp(31552) := x"21e3";
    tmp(31553) := x"2a03";
    tmp(31554) := x"2a03";
    tmp(31555) := x"21e2";
    tmp(31556) := x"1181";
    tmp(31557) := x"1141";
    tmp(31558) := x"1121";
    tmp(31559) := x"1121";
    tmp(31560) := x"1141";
    tmp(31561) := x"1121";
    tmp(31562) := x"1141";
    tmp(31563) := x"1120";
    tmp(31564) := x"1100";
    tmp(31565) := x"1120";
    tmp(31566) := x"1120";
    tmp(31567) := x"1141";
    tmp(31568) := x"1141";
    tmp(31569) := x"1961";
    tmp(31570) := x"1982";
    tmp(31571) := x"1981";
    tmp(31572) := x"1941";
    tmp(31573) := x"1941";
    tmp(31574) := x"1121";
    tmp(31575) := x"1120";
    tmp(31576) := x"1120";
    tmp(31577) := x"1921";
    tmp(31578) := x"1921";
    tmp(31579) := x"1941";
    tmp(31580) := x"2161";
    tmp(31581) := x"2181";
    tmp(31582) := x"29a2";
    tmp(31583) := x"31c2";
    tmp(31584) := x"39e2";
    tmp(31585) := x"39e3";
    tmp(31586) := x"39e3";
    tmp(31587) := x"31c2";
    tmp(31588) := x"31c3";
    tmp(31589) := x"39c3";
    tmp(31590) := x"31a3";
    tmp(31591) := x"3182";
    tmp(31592) := x"2962";
    tmp(31593) := x"2962";
    tmp(31594) := x"2962";
    tmp(31595) := x"2942";
    tmp(31596) := x"2142";
    tmp(31597) := x"2942";
    tmp(31598) := x"2962";
    tmp(31599) := x"2962";
    tmp(31600) := x"2963";
    tmp(31601) := x"2962";
    tmp(31602) := x"2962";
    tmp(31603) := x"2962";
    tmp(31604) := x"3163";
    tmp(31605) := x"2963";
    tmp(31606) := x"2963";
    tmp(31607) := x"2963";
    tmp(31608) := x"2942";
    tmp(31609) := x"2122";
    tmp(31610) := x"2102";
    tmp(31611) := x"2102";
    tmp(31612) := x"2903";
    tmp(31613) := x"2903";
    tmp(31614) := x"2903";
    tmp(31615) := x"2923";
    tmp(31616) := x"2923";
    tmp(31617) := x"2923";
    tmp(31618) := x"3124";
    tmp(31619) := x"3144";
    tmp(31620) := x"3144";
    tmp(31621) := x"3944";
    tmp(31622) := x"3945";
    tmp(31623) := x"3944";
    tmp(31624) := x"3965";
    tmp(31625) := x"3965";
    tmp(31626) := x"3985";
    tmp(31627) := x"4186";
    tmp(31628) := x"41a6";
    tmp(31629) := x"41a7";
    tmp(31630) := x"49c7";
    tmp(31631) := x"49e7";
    tmp(31632) := x"49e7";
    tmp(31633) := x"5208";
    tmp(31634) := x"5208";
    tmp(31635) := x"5209";
    tmp(31636) := x"5229";
    tmp(31637) := x"07e0";
    tmp(31638) := x"07e0";
    tmp(31639) := x"07e0";
    tmp(31640) := x"07e0";
    tmp(31641) := x"07e0";
    tmp(31642) := x"07e0";
    tmp(31643) := x"07e0";
    tmp(31644) := x"07e0";
    tmp(31645) := x"07e0";
    tmp(31646) := x"07e0";
    tmp(31647) := x"07e0";
    tmp(31648) := x"07e0";
    tmp(31649) := x"07e0";
    tmp(31650) := x"07e0";
    tmp(31651) := x"07e0";
    tmp(31652) := x"07e0";
    tmp(31653) := x"07e0";
    tmp(31654) := x"07e0";
    tmp(31655) := x"07e0";
    tmp(31656) := x"07e0";
    tmp(31657) := x"07e0";
    tmp(31658) := x"07e0";
    tmp(31659) := x"07e0";
    tmp(31660) := x"07e0";
    tmp(31661) := x"07e0";
    tmp(31662) := x"07e0";
    tmp(31663) := x"07e0";
    tmp(31664) := x"07e0";
    tmp(31665) := x"07e0";
    tmp(31666) := x"07e0";
    tmp(31667) := x"07e0";
    tmp(31668) := x"07e0";
    tmp(31669) := x"07e0";
    tmp(31670) := x"07e0";
    tmp(31671) := x"07e0";
    tmp(31672) := x"07e0";
    tmp(31673) := x"07e0";
    tmp(31674) := x"07e0";
    tmp(31675) := x"07e0";
    tmp(31676) := x"07e0";
    tmp(31677) := x"0840";
    tmp(31678) := x"0840";
    tmp(31679) := x"0840";
    tmp(31680) := x"0000";
    tmp(31681) := x"00c5";
    tmp(31682) := x"00e5";
    tmp(31683) := x"00e5";
    tmp(31684) := x"00e5";
    tmp(31685) := x"00c5";
    tmp(31686) := x"00c4";
    tmp(31687) := x"00a4";
    tmp(31688) := x"00a4";
    tmp(31689) := x"0083";
    tmp(31690) := x"0082";
    tmp(31691) := x"0082";
    tmp(31692) := x"00a3";
    tmp(31693) := x"00a3";
    tmp(31694) := x"0062";
    tmp(31695) := x"0041";
    tmp(31696) := x"0021";
    tmp(31697) := x"0041";
    tmp(31698) := x"0882";
    tmp(31699) := x"0062";
    tmp(31700) := x"0062";
    tmp(31701) := x"0862";
    tmp(31702) := x"0882";
    tmp(31703) := x"0062";
    tmp(31704) := x"08a3";
    tmp(31705) := x"0926";
    tmp(31706) := x"0905";
    tmp(31707) := x"0905";
    tmp(31708) := x"0905";
    tmp(31709) := x"0905";
    tmp(31710) := x"08e4";
    tmp(31711) := x"08e4";
    tmp(31712) := x"08e5";
    tmp(31713) := x"0905";
    tmp(31714) := x"0905";
    tmp(31715) := x"0926";
    tmp(31716) := x"0905";
    tmp(31717) := x"08e4";
    tmp(31718) := x"08c4";
    tmp(31719) := x"08c4";
    tmp(31720) := x"0905";
    tmp(31721) := x"0926";
    tmp(31722) := x"0925";
    tmp(31723) := x"0925";
    tmp(31724) := x"0925";
    tmp(31725) := x"0904";
    tmp(31726) := x"08e4";
    tmp(31727) := x"08c3";
    tmp(31728) := x"08c3";
    tmp(31729) := x"08e4";
    tmp(31730) := x"0925";
    tmp(31731) := x"0904";
    tmp(31732) := x"08e4";
    tmp(31733) := x"08e3";
    tmp(31734) := x"08e3";
    tmp(31735) := x"1104";
    tmp(31736) := x"08a2";
    tmp(31737) := x"08c2";
    tmp(31738) := x"1142";
    tmp(31739) := x"1121";
    tmp(31740) := x"1120";
    tmp(31741) := x"1120";
    tmp(31742) := x"0920";
    tmp(31743) := x"0920";
    tmp(31744) := x"0900";
    tmp(31745) := x"0920";
    tmp(31746) := x"0900";
    tmp(31747) := x"0920";
    tmp(31748) := x"0900";
    tmp(31749) := x"0900";
    tmp(31750) := x"0900";
    tmp(31751) := x"08e0";
    tmp(31752) := x"0900";
    tmp(31753) := x"1101";
    tmp(31754) := x"1121";
    tmp(31755) := x"1962";
    tmp(31756) := x"2183";
    tmp(31757) := x"21a3";
    tmp(31758) := x"31e4";
    tmp(31759) := x"3226";
    tmp(31760) := x"3a26";
    tmp(31761) := x"4248";
    tmp(31762) := x"4a89";
    tmp(31763) := x"52aa";
    tmp(31764) := x"5acb";
    tmp(31765) := x"5aab";
    tmp(31766) := x"5acb";
    tmp(31767) := x"5aec";
    tmp(31768) := x"62ed";
    tmp(31769) := x"6b2f";
    tmp(31770) := x"6b2f";
    tmp(31771) := x"632e";
    tmp(31772) := x"6b2f";
    tmp(31773) := x"630f";
    tmp(31774) := x"5aee";
    tmp(31775) := x"5acd";
    tmp(31776) := x"5acb";
    tmp(31777) := x"52a9";
    tmp(31778) := x"5288";
    tmp(31779) := x"4a87";
    tmp(31780) := x"4226";
    tmp(31781) := x"39e5";
    tmp(31782) := x"31c4";
    tmp(31783) := x"2983";
    tmp(31784) := x"21a3";
    tmp(31785) := x"2183";
    tmp(31786) := x"2184";
    tmp(31787) := x"21a4";
    tmp(31788) := x"19a4";
    tmp(31789) := x"1984";
    tmp(31790) := x"19a3";
    tmp(31791) := x"21a3";
    tmp(31792) := x"29e3";
    tmp(31793) := x"29e3";
    tmp(31794) := x"21e2";
    tmp(31795) := x"19a1";
    tmp(31796) := x"1141";
    tmp(31797) := x"1141";
    tmp(31798) := x"1141";
    tmp(31799) := x"1121";
    tmp(31800) := x"1121";
    tmp(31801) := x"1141";
    tmp(31802) := x"1121";
    tmp(31803) := x"1120";
    tmp(31804) := x"1100";
    tmp(31805) := x"1100";
    tmp(31806) := x"1120";
    tmp(31807) := x"1120";
    tmp(31808) := x"1141";
    tmp(31809) := x"1941";
    tmp(31810) := x"1961";
    tmp(31811) := x"1961";
    tmp(31812) := x"1961";
    tmp(31813) := x"1941";
    tmp(31814) := x"1121";
    tmp(31815) := x"1120";
    tmp(31816) := x"1120";
    tmp(31817) := x"1120";
    tmp(31818) := x"1941";
    tmp(31819) := x"1941";
    tmp(31820) := x"1941";
    tmp(31821) := x"2141";
    tmp(31822) := x"2161";
    tmp(31823) := x"2981";
    tmp(31824) := x"29a2";
    tmp(31825) := x"31a2";
    tmp(31826) := x"31a2";
    tmp(31827) := x"31a2";
    tmp(31828) := x"31a2";
    tmp(31829) := x"3182";
    tmp(31830) := x"3183";
    tmp(31831) := x"2982";
    tmp(31832) := x"2942";
    tmp(31833) := x"2942";
    tmp(31834) := x"2942";
    tmp(31835) := x"2942";
    tmp(31836) := x"2142";
    tmp(31837) := x"2142";
    tmp(31838) := x"2942";
    tmp(31839) := x"2962";
    tmp(31840) := x"2942";
    tmp(31841) := x"2963";
    tmp(31842) := x"2963";
    tmp(31843) := x"2963";
    tmp(31844) := x"3163";
    tmp(31845) := x"2963";
    tmp(31846) := x"2942";
    tmp(31847) := x"2943";
    tmp(31848) := x"2942";
    tmp(31849) := x"2122";
    tmp(31850) := x"2102";
    tmp(31851) := x"2102";
    tmp(31852) := x"2103";
    tmp(31853) := x"2903";
    tmp(31854) := x"2903";
    tmp(31855) := x"2903";
    tmp(31856) := x"2903";
    tmp(31857) := x"2923";
    tmp(31858) := x"3123";
    tmp(31859) := x"3123";
    tmp(31860) := x"3124";
    tmp(31861) := x"3123";
    tmp(31862) := x"3124";
    tmp(31863) := x"3124";
    tmp(31864) := x"3124";
    tmp(31865) := x"3124";
    tmp(31866) := x"3124";
    tmp(31867) := x"3144";
    tmp(31868) := x"3144";
    tmp(31869) := x"3144";
    tmp(31870) := x"3965";
    tmp(31871) := x"3965";
    tmp(31872) := x"3985";
    tmp(31873) := x"4186";
    tmp(31874) := x"4186";
    tmp(31875) := x"41c6";
    tmp(31876) := x"41a6";
    tmp(31877) := x"07e0";
    tmp(31878) := x"07e0";
    tmp(31879) := x"07e0";
    tmp(31880) := x"07e0";
    tmp(31881) := x"07e0";
    tmp(31882) := x"07e0";
    tmp(31883) := x"07e0";
    tmp(31884) := x"07e0";
    tmp(31885) := x"07e0";
    tmp(31886) := x"07e0";
    tmp(31887) := x"07e0";
    tmp(31888) := x"07e0";
    tmp(31889) := x"07e0";
    tmp(31890) := x"07e0";
    tmp(31891) := x"07e0";
    tmp(31892) := x"07e0";
    tmp(31893) := x"07e0";
    tmp(31894) := x"07e0";
    tmp(31895) := x"07e0";
    tmp(31896) := x"07e0";
    tmp(31897) := x"07e0";
    tmp(31898) := x"07e0";
    tmp(31899) := x"07e0";
    tmp(31900) := x"07e0";
    tmp(31901) := x"07e0";
    tmp(31902) := x"07e0";
    tmp(31903) := x"07e0";
    tmp(31904) := x"07e0";
    tmp(31905) := x"07e0";
    tmp(31906) := x"07e0";
    tmp(31907) := x"07e0";
    tmp(31908) := x"07e0";
    tmp(31909) := x"07e0";
    tmp(31910) := x"07e0";
    tmp(31911) := x"07e0";
    tmp(31912) := x"07e0";
    tmp(31913) := x"07e0";
    tmp(31914) := x"07e0";
    tmp(31915) := x"07e0";
    tmp(31916) := x"07e0";
    tmp(31917) := x"0840";
    tmp(31918) := x"0840";
    tmp(31919) := x"0840";
    tmp(31920) := x"0020";
    tmp(31921) := x"00c4";
    tmp(31922) := x"00a4";
    tmp(31923) := x"00c5";
    tmp(31924) := x"0106";
    tmp(31925) := x"0106";
    tmp(31926) := x"00e5";
    tmp(31927) := x"00e5";
    tmp(31928) := x"00c5";
    tmp(31929) := x"00a3";
    tmp(31930) := x"0083";
    tmp(31931) := x"00a3";
    tmp(31932) := x"00a4";
    tmp(31933) := x"00a4";
    tmp(31934) := x"00c4";
    tmp(31935) := x"00c4";
    tmp(31936) := x"00a3";
    tmp(31937) := x"0062";
    tmp(31938) := x"0062";
    tmp(31939) := x"0041";
    tmp(31940) := x"0041";
    tmp(31941) := x"0021";
    tmp(31942) := x"0041";
    tmp(31943) := x"0082";
    tmp(31944) := x"0905";
    tmp(31945) := x"0925";
    tmp(31946) := x"0905";
    tmp(31947) := x"0905";
    tmp(31948) := x"0926";
    tmp(31949) := x"0926";
    tmp(31950) := x"0926";
    tmp(31951) := x"08e5";
    tmp(31952) := x"00c4";
    tmp(31953) := x"0905";
    tmp(31954) := x"0905";
    tmp(31955) := x"0905";
    tmp(31956) := x"08e4";
    tmp(31957) := x"08e4";
    tmp(31958) := x"08e4";
    tmp(31959) := x"0905";
    tmp(31960) := x"0926";
    tmp(31961) := x"0946";
    tmp(31962) := x"0925";
    tmp(31963) := x"0925";
    tmp(31964) := x"0925";
    tmp(31965) := x"0924";
    tmp(31966) := x"0904";
    tmp(31967) := x"08e3";
    tmp(31968) := x"08c3";
    tmp(31969) := x"0904";
    tmp(31970) := x"0925";
    tmp(31971) := x"1145";
    tmp(31972) := x"0924";
    tmp(31973) := x"08e3";
    tmp(31974) := x"08e3";
    tmp(31975) := x"08a2";
    tmp(31976) := x"08a2";
    tmp(31977) := x"1102";
    tmp(31978) := x"1121";
    tmp(31979) := x"1120";
    tmp(31980) := x"1120";
    tmp(31981) := x"1120";
    tmp(31982) := x"1120";
    tmp(31983) := x"0920";
    tmp(31984) := x"1120";
    tmp(31985) := x"1120";
    tmp(31986) := x"0920";
    tmp(31987) := x"0920";
    tmp(31988) := x"0900";
    tmp(31989) := x"0900";
    tmp(31990) := x"0900";
    tmp(31991) := x"08e0";
    tmp(31992) := x"08e0";
    tmp(31993) := x"0900";
    tmp(31994) := x"1121";
    tmp(31995) := x"1141";
    tmp(31996) := x"1942";
    tmp(31997) := x"2183";
    tmp(31998) := x"29a4";
    tmp(31999) := x"29c4";
    tmp(32000) := x"31c5";
    tmp(32001) := x"3a26";
    tmp(32002) := x"4247";
    tmp(32003) := x"4a48";
    tmp(32004) := x"4a69";
    tmp(32005) := x"5269";
    tmp(32006) := x"528a";
    tmp(32007) := x"528b";
    tmp(32008) := x"5acd";
    tmp(32009) := x"62cd";
    tmp(32010) := x"5acd";
    tmp(32011) := x"5acd";
    tmp(32012) := x"5acd";
    tmp(32013) := x"5acc";
    tmp(32014) := x"5aac";
    tmp(32015) := x"528b";
    tmp(32016) := x"5289";
    tmp(32017) := x"4a88";
    tmp(32018) := x"4a67";
    tmp(32019) := x"4206";
    tmp(32020) := x"39e5";
    tmp(32021) := x"31c4";
    tmp(32022) := x"29a4";
    tmp(32023) := x"2984";
    tmp(32024) := x"2184";
    tmp(32025) := x"2184";
    tmp(32026) := x"21a4";
    tmp(32027) := x"21c5";
    tmp(32028) := x"21a4";
    tmp(32029) := x"1983";
    tmp(32030) := x"1983";
    tmp(32031) := x"21c3";
    tmp(32032) := x"21e3";
    tmp(32033) := x"21c2";
    tmp(32034) := x"21a1";
    tmp(32035) := x"1141";
    tmp(32036) := x"1121";
    tmp(32037) := x"1121";
    tmp(32038) := x"1141";
    tmp(32039) := x"1121";
    tmp(32040) := x"1121";
    tmp(32041) := x"1121";
    tmp(32042) := x"1121";
    tmp(32043) := x"1120";
    tmp(32044) := x"1120";
    tmp(32045) := x"1100";
    tmp(32046) := x"1120";
    tmp(32047) := x"1120";
    tmp(32048) := x"1120";
    tmp(32049) := x"1141";
    tmp(32050) := x"1961";
    tmp(32051) := x"1961";
    tmp(32052) := x"1961";
    tmp(32053) := x"1941";
    tmp(32054) := x"1921";
    tmp(32055) := x"1121";
    tmp(32056) := x"1120";
    tmp(32057) := x"1120";
    tmp(32058) := x"1920";
    tmp(32059) := x"1941";
    tmp(32060) := x"1941";
    tmp(32061) := x"1941";
    tmp(32062) := x"2141";
    tmp(32063) := x"2161";
    tmp(32064) := x"2981";
    tmp(32065) := x"2982";
    tmp(32066) := x"2982";
    tmp(32067) := x"2982";
    tmp(32068) := x"2982";
    tmp(32069) := x"2962";
    tmp(32070) := x"2982";
    tmp(32071) := x"2962";
    tmp(32072) := x"2142";
    tmp(32073) := x"2121";
    tmp(32074) := x"2101";
    tmp(32075) := x"2121";
    tmp(32076) := x"2121";
    tmp(32077) := x"2122";
    tmp(32078) := x"2142";
    tmp(32079) := x"2142";
    tmp(32080) := x"2962";
    tmp(32081) := x"2963";
    tmp(32082) := x"2983";
    tmp(32083) := x"2963";
    tmp(32084) := x"2963";
    tmp(32085) := x"2962";
    tmp(32086) := x"2942";
    tmp(32087) := x"2942";
    tmp(32088) := x"2122";
    tmp(32089) := x"2122";
    tmp(32090) := x"2102";
    tmp(32091) := x"2102";
    tmp(32092) := x"2903";
    tmp(32093) := x"2903";
    tmp(32094) := x"2903";
    tmp(32095) := x"2903";
    tmp(32096) := x"2903";
    tmp(32097) := x"2903";
    tmp(32098) := x"2903";
    tmp(32099) := x"2903";
    tmp(32100) := x"2903";
    tmp(32101) := x"2903";
    tmp(32102) := x"28e3";
    tmp(32103) := x"28e3";
    tmp(32104) := x"28e3";
    tmp(32105) := x"28e3";
    tmp(32106) := x"28e3";
    tmp(32107) := x"28e3";
    tmp(32108) := x"28e3";
    tmp(32109) := x"2903";
    tmp(32110) := x"2903";
    tmp(32111) := x"2903";
    tmp(32112) := x"3124";
    tmp(32113) := x"3124";
    tmp(32114) := x"3124";
    tmp(32115) := x"3944";
    tmp(32116) := x"3945";
    tmp(32117) := x"07e0";
    tmp(32118) := x"07e0";
    tmp(32119) := x"07e0";
    tmp(32120) := x"07e0";
    tmp(32121) := x"07e0";
    tmp(32122) := x"07e0";
    tmp(32123) := x"07e0";
    tmp(32124) := x"07e0";
    tmp(32125) := x"07e0";
    tmp(32126) := x"07e0";
    tmp(32127) := x"07e0";
    tmp(32128) := x"07e0";
    tmp(32129) := x"07e0";
    tmp(32130) := x"07e0";
    tmp(32131) := x"07e0";
    tmp(32132) := x"07e0";
    tmp(32133) := x"07e0";
    tmp(32134) := x"07e0";
    tmp(32135) := x"07e0";
    tmp(32136) := x"07e0";
    tmp(32137) := x"07e0";
    tmp(32138) := x"07e0";
    tmp(32139) := x"07e0";
    tmp(32140) := x"07e0";
    tmp(32141) := x"07e0";
    tmp(32142) := x"07e0";
    tmp(32143) := x"07e0";
    tmp(32144) := x"07e0";
    tmp(32145) := x"07e0";
    tmp(32146) := x"07e0";
    tmp(32147) := x"07e0";
    tmp(32148) := x"07e0";
    tmp(32149) := x"07e0";
    tmp(32150) := x"07e0";
    tmp(32151) := x"07e0";
    tmp(32152) := x"07e0";
    tmp(32153) := x"07e0";
    tmp(32154) := x"07e0";
    tmp(32155) := x"07e0";
    tmp(32156) := x"07e0";
    tmp(32157) := x"0840";
    tmp(32158) := x"0840";
    tmp(32159) := x"0840";
    tmp(32160) := x"0020";
    tmp(32161) := x"00e5";
    tmp(32162) := x"00e5";
    tmp(32163) := x"00c5";
    tmp(32164) := x"00c4";
    tmp(32165) := x"00c5";
    tmp(32166) := x"00e5";
    tmp(32167) := x"00e5";
    tmp(32168) := x"00e5";
    tmp(32169) := x"00e5";
    tmp(32170) := x"00a4";
    tmp(32171) := x"00a4";
    tmp(32172) := x"00a4";
    tmp(32173) := x"00c4";
    tmp(32174) := x"00c4";
    tmp(32175) := x"00e5";
    tmp(32176) := x"00c4";
    tmp(32177) := x"00c4";
    tmp(32178) := x"00c4";
    tmp(32179) := x"08a3";
    tmp(32180) := x"0082";
    tmp(32181) := x"0062";
    tmp(32182) := x"0082";
    tmp(32183) := x"08e4";
    tmp(32184) := x"0926";
    tmp(32185) := x"0946";
    tmp(32186) := x"0906";
    tmp(32187) := x"0905";
    tmp(32188) := x"0905";
    tmp(32189) := x"0905";
    tmp(32190) := x"08e4";
    tmp(32191) := x"00c4";
    tmp(32192) := x"08e5";
    tmp(32193) := x"08e5";
    tmp(32194) := x"08e5";
    tmp(32195) := x"0905";
    tmp(32196) := x"0905";
    tmp(32197) := x"0905";
    tmp(32198) := x"0905";
    tmp(32199) := x"0905";
    tmp(32200) := x"0925";
    tmp(32201) := x"0946";
    tmp(32202) := x"0925";
    tmp(32203) := x"0925";
    tmp(32204) := x"0925";
    tmp(32205) := x"0904";
    tmp(32206) := x"0904";
    tmp(32207) := x"08e4";
    tmp(32208) := x"0904";
    tmp(32209) := x"0904";
    tmp(32210) := x"0925";
    tmp(32211) := x"0904";
    tmp(32212) := x"0904";
    tmp(32213) := x"0924";
    tmp(32214) := x"1124";
    tmp(32215) := x"08c2";
    tmp(32216) := x"1102";
    tmp(32217) := x"1121";
    tmp(32218) := x"1141";
    tmp(32219) := x"1140";
    tmp(32220) := x"1140";
    tmp(32221) := x"1120";
    tmp(32222) := x"1120";
    tmp(32223) := x"1120";
    tmp(32224) := x"1120";
    tmp(32225) := x"1120";
    tmp(32226) := x"0920";
    tmp(32227) := x"0920";
    tmp(32228) := x"0900";
    tmp(32229) := x"0900";
    tmp(32230) := x"0900";
    tmp(32231) := x"0900";
    tmp(32232) := x"08e0";
    tmp(32233) := x"0900";
    tmp(32234) := x"1121";
    tmp(32235) := x"1121";
    tmp(32236) := x"1122";
    tmp(32237) := x"1962";
    tmp(32238) := x"2183";
    tmp(32239) := x"29a4";
    tmp(32240) := x"31c4";
    tmp(32241) := x"31e5";
    tmp(32242) := x"3a06";
    tmp(32243) := x"3a06";
    tmp(32244) := x"4227";
    tmp(32245) := x"4a48";
    tmp(32246) := x"4a68";
    tmp(32247) := x"528a";
    tmp(32248) := x"528a";
    tmp(32249) := x"528b";
    tmp(32250) := x"528b";
    tmp(32251) := x"528c";
    tmp(32252) := x"528b";
    tmp(32253) := x"528a";
    tmp(32254) := x"526a";
    tmp(32255) := x"4a49";
    tmp(32256) := x"4a48";
    tmp(32257) := x"4227";
    tmp(32258) := x"3a06";
    tmp(32259) := x"31c5";
    tmp(32260) := x"31c5";
    tmp(32261) := x"29a4";
    tmp(32262) := x"2984";
    tmp(32263) := x"29a4";
    tmp(32264) := x"21a4";
    tmp(32265) := x"21a4";
    tmp(32266) := x"29e5";
    tmp(32267) := x"21c5";
    tmp(32268) := x"1984";
    tmp(32269) := x"1983";
    tmp(32270) := x"21a3";
    tmp(32271) := x"21c3";
    tmp(32272) := x"21c2";
    tmp(32273) := x"21a2";
    tmp(32274) := x"1961";
    tmp(32275) := x"1121";
    tmp(32276) := x"1121";
    tmp(32277) := x"1121";
    tmp(32278) := x"1141";
    tmp(32279) := x"1121";
    tmp(32280) := x"1120";
    tmp(32281) := x"1120";
    tmp(32282) := x"1120";
    tmp(32283) := x"1120";
    tmp(32284) := x"1120";
    tmp(32285) := x"1100";
    tmp(32286) := x"1100";
    tmp(32287) := x"1120";
    tmp(32288) := x"1120";
    tmp(32289) := x"1120";
    tmp(32290) := x"1141";
    tmp(32291) := x"1961";
    tmp(32292) := x"1961";
    tmp(32293) := x"1941";
    tmp(32294) := x"1941";
    tmp(32295) := x"1121";
    tmp(32296) := x"1120";
    tmp(32297) := x"1120";
    tmp(32298) := x"1120";
    tmp(32299) := x"1940";
    tmp(32300) := x"1940";
    tmp(32301) := x"1921";
    tmp(32302) := x"1941";
    tmp(32303) := x"1941";
    tmp(32304) := x"2141";
    tmp(32305) := x"2161";
    tmp(32306) := x"2161";
    tmp(32307) := x"2961";
    tmp(32308) := x"2141";
    tmp(32309) := x"2142";
    tmp(32310) := x"2962";
    tmp(32311) := x"2142";
    tmp(32312) := x"2122";
    tmp(32313) := x"1901";
    tmp(32314) := x"18e1";
    tmp(32315) := x"18e1";
    tmp(32316) := x"1901";
    tmp(32317) := x"2101";
    tmp(32318) := x"2122";
    tmp(32319) := x"2142";
    tmp(32320) := x"2962";
    tmp(32321) := x"2962";
    tmp(32322) := x"2963";
    tmp(32323) := x"2963";
    tmp(32324) := x"2962";
    tmp(32325) := x"2942";
    tmp(32326) := x"2922";
    tmp(32327) := x"2922";
    tmp(32328) := x"2122";
    tmp(32329) := x"2102";
    tmp(32330) := x"2102";
    tmp(32331) := x"2102";
    tmp(32332) := x"2903";
    tmp(32333) := x"2903";
    tmp(32334) := x"2102";
    tmp(32335) := x"20e3";
    tmp(32336) := x"20e2";
    tmp(32337) := x"20e2";
    tmp(32338) := x"20e2";
    tmp(32339) := x"20e2";
    tmp(32340) := x"28e2";
    tmp(32341) := x"20c2";
    tmp(32342) := x"20c2";
    tmp(32343) := x"20c2";
    tmp(32344) := x"20c2";
    tmp(32345) := x"20c2";
    tmp(32346) := x"20c2";
    tmp(32347) := x"20c2";
    tmp(32348) := x"20a2";
    tmp(32349) := x"20c2";
    tmp(32350) := x"20c2";
    tmp(32351) := x"20e2";
    tmp(32352) := x"20e2";
    tmp(32353) := x"28e3";
    tmp(32354) := x"28e3";
    tmp(32355) := x"2903";
    tmp(32356) := x"2903";
    tmp(32357) := x"07e0";
    tmp(32358) := x"07e0";
    tmp(32359) := x"07e0";
    tmp(32360) := x"07e0";
    tmp(32361) := x"07e0";
    tmp(32362) := x"07e0";
    tmp(32363) := x"07e0";
    tmp(32364) := x"07e0";
    tmp(32365) := x"07e0";
    tmp(32366) := x"07e0";
    tmp(32367) := x"07e0";
    tmp(32368) := x"07e0";
    tmp(32369) := x"07e0";
    tmp(32370) := x"07e0";
    tmp(32371) := x"07e0";
    tmp(32372) := x"07e0";
    tmp(32373) := x"07e0";
    tmp(32374) := x"07e0";
    tmp(32375) := x"07e0";
    tmp(32376) := x"07e0";
    tmp(32377) := x"07e0";
    tmp(32378) := x"07e0";
    tmp(32379) := x"07e0";
    tmp(32380) := x"07e0";
    tmp(32381) := x"07e0";
    tmp(32382) := x"07e0";
    tmp(32383) := x"07e0";
    tmp(32384) := x"07e0";
    tmp(32385) := x"07e0";
    tmp(32386) := x"07e0";
    tmp(32387) := x"07e0";
    tmp(32388) := x"07e0";
    tmp(32389) := x"07e0";
    tmp(32390) := x"07e0";
    tmp(32391) := x"07e0";
    tmp(32392) := x"07e0";
    tmp(32393) := x"07e0";
    tmp(32394) := x"07e0";
    tmp(32395) := x"07e0";
    tmp(32396) := x"07e0";
    tmp(32397) := x"0840";
    tmp(32398) := x"0840";
    tmp(32399) := x"0840";
    tmp(32400) := x"0020";
    tmp(32401) := x"00e5";
    tmp(32402) := x"00e5";
    tmp(32403) := x"00c4";
    tmp(32404) := x"00c5";
    tmp(32405) := x"00c5";
    tmp(32406) := x"00c5";
    tmp(32407) := x"00e5";
    tmp(32408) := x"00e6";
    tmp(32409) := x"0106";
    tmp(32410) := x"00e5";
    tmp(32411) := x"00c5";
    tmp(32412) := x"00c5";
    tmp(32413) := x"00e5";
    tmp(32414) := x"00e5";
    tmp(32415) := x"0105";
    tmp(32416) := x"00e5";
    tmp(32417) := x"00e5";
    tmp(32418) := x"00c5";
    tmp(32419) := x"00e5";
    tmp(32420) := x"0905";
    tmp(32421) := x"08e5";
    tmp(32422) := x"08e5";
    tmp(32423) := x"08e5";
    tmp(32424) := x"0905";
    tmp(32425) := x"0905";
    tmp(32426) := x"08e5";
    tmp(32427) := x"08e4";
    tmp(32428) := x"08e4";
    tmp(32429) := x"08e4";
    tmp(32430) := x"08c4";
    tmp(32431) := x"08e5";
    tmp(32432) := x"0905";
    tmp(32433) := x"0905";
    tmp(32434) := x"0905";
    tmp(32435) := x"0905";
    tmp(32436) := x"0905";
    tmp(32437) := x"0925";
    tmp(32438) := x"0905";
    tmp(32439) := x"0905";
    tmp(32440) := x"0905";
    tmp(32441) := x"0925";
    tmp(32442) := x"0925";
    tmp(32443) := x"0925";
    tmp(32444) := x"0925";
    tmp(32445) := x"0905";
    tmp(32446) := x"0904";
    tmp(32447) := x"0925";
    tmp(32448) := x"0905";
    tmp(32449) := x"0904";
    tmp(32450) := x"0925";
    tmp(32451) := x"0904";
    tmp(32452) := x"08c3";
    tmp(32453) := x"08e3";
    tmp(32454) := x"08c2";
    tmp(32455) := x"08e1";
    tmp(32456) := x"1141";
    tmp(32457) := x"1141";
    tmp(32458) := x"1141";
    tmp(32459) := x"1140";
    tmp(32460) := x"1140";
    tmp(32461) := x"1120";
    tmp(32462) := x"1120";
    tmp(32463) := x"1120";
    tmp(32464) := x"1120";
    tmp(32465) := x"1120";
    tmp(32466) := x"1120";
    tmp(32467) := x"1120";
    tmp(32468) := x"0920";
    tmp(32469) := x"0900";
    tmp(32470) := x"0900";
    tmp(32471) := x"0900";
    tmp(32472) := x"0900";
    tmp(32473) := x"08e0";
    tmp(32474) := x"1101";
    tmp(32475) := x"1101";
    tmp(32476) := x"1121";
    tmp(32477) := x"1922";
    tmp(32478) := x"1962";
    tmp(32479) := x"2183";
    tmp(32480) := x"29a3";
    tmp(32481) := x"29a4";
    tmp(32482) := x"31a5";
    tmp(32483) := x"31e5";
    tmp(32484) := x"39e6";
    tmp(32485) := x"4227";
    tmp(32486) := x"4248";
    tmp(32487) := x"4a48";
    tmp(32488) := x"4a49";
    tmp(32489) := x"4a49";
    tmp(32490) := x"4a6a";
    tmp(32491) := x"4a4a";
    tmp(32492) := x"4a49";
    tmp(32493) := x"4a48";
    tmp(32494) := x"4228";
    tmp(32495) := x"4207";
    tmp(32496) := x"3a06";
    tmp(32497) := x"3a06";
    tmp(32498) := x"31c5";
    tmp(32499) := x"31a5";
    tmp(32500) := x"29a5";
    tmp(32501) := x"2985";
    tmp(32502) := x"2984";
    tmp(32503) := x"29a5";
    tmp(32504) := x"29c5";
    tmp(32505) := x"29e5";
    tmp(32506) := x"29e5";
    tmp(32507) := x"21a4";
    tmp(32508) := x"1963";
    tmp(32509) := x"1983";
    tmp(32510) := x"21a3";
    tmp(32511) := x"21c2";
    tmp(32512) := x"1982";
    tmp(32513) := x"1961";
    tmp(32514) := x"1121";
    tmp(32515) := x"1121";
    tmp(32516) := x"1121";
    tmp(32517) := x"1121";
    tmp(32518) := x"1121";
    tmp(32519) := x"1120";
    tmp(32520) := x"1120";
    tmp(32521) := x"1100";
    tmp(32522) := x"1120";
    tmp(32523) := x"1120";
    tmp(32524) := x"1120";
    tmp(32525) := x"1100";
    tmp(32526) := x"1100";
    tmp(32527) := x"1100";
    tmp(32528) := x"1100";
    tmp(32529) := x"1120";
    tmp(32530) := x"1140";
    tmp(32531) := x"1141";
    tmp(32532) := x"1141";
    tmp(32533) := x"1141";
    tmp(32534) := x"1941";
    tmp(32535) := x"1121";
    tmp(32536) := x"1120";
    tmp(32537) := x"1120";
    tmp(32538) := x"1120";
    tmp(32539) := x"1920";
    tmp(32540) := x"1940";
    tmp(32541) := x"1921";
    tmp(32542) := x"1921";
    tmp(32543) := x"1921";
    tmp(32544) := x"2121";
    tmp(32545) := x"2141";
    tmp(32546) := x"2141";
    tmp(32547) := x"2141";
    tmp(32548) := x"2141";
    tmp(32549) := x"2141";
    tmp(32550) := x"2121";
    tmp(32551) := x"2142";
    tmp(32552) := x"2121";
    tmp(32553) := x"18e1";
    tmp(32554) := x"18c1";
    tmp(32555) := x"18c1";
    tmp(32556) := x"18e1";
    tmp(32557) := x"1901";
    tmp(32558) := x"2122";
    tmp(32559) := x"2142";
    tmp(32560) := x"2942";
    tmp(32561) := x"2962";
    tmp(32562) := x"2962";
    tmp(32563) := x"2942";
    tmp(32564) := x"2142";
    tmp(32565) := x"2122";
    tmp(32566) := x"2122";
    tmp(32567) := x"2122";
    tmp(32568) := x"2122";
    tmp(32569) := x"2102";
    tmp(32570) := x"2122";
    tmp(32571) := x"2102";
    tmp(32572) := x"2102";
    tmp(32573) := x"20e2";
    tmp(32574) := x"20e2";
    tmp(32575) := x"20e2";
    tmp(32576) := x"20c2";
    tmp(32577) := x"20c2";
    tmp(32578) := x"20c2";
    tmp(32579) := x"20c2";
    tmp(32580) := x"20c2";
    tmp(32581) := x"20a2";
    tmp(32582) := x"20a2";
    tmp(32583) := x"18a2";
    tmp(32584) := x"18a1";
    tmp(32585) := x"18a1";
    tmp(32586) := x"18a1";
    tmp(32587) := x"18a1";
    tmp(32588) := x"18a1";
    tmp(32589) := x"18a1";
    tmp(32590) := x"18a1";
    tmp(32591) := x"20a2";
    tmp(32592) := x"20c2";
    tmp(32593) := x"20c2";
    tmp(32594) := x"20c2";
    tmp(32595) := x"20e2";
    tmp(32596) := x"20e2";
    tmp(32597) := x"07e0";
    tmp(32598) := x"07e0";
    tmp(32599) := x"07e0";
    tmp(32600) := x"07e0";
    tmp(32601) := x"07e0";
    tmp(32602) := x"07e0";
    tmp(32603) := x"07e0";
    tmp(32604) := x"07e0";
    tmp(32605) := x"07e0";
    tmp(32606) := x"07e0";
    tmp(32607) := x"07e0";
    tmp(32608) := x"07e0";
    tmp(32609) := x"07e0";
    tmp(32610) := x"07e0";
    tmp(32611) := x"07e0";
    tmp(32612) := x"07e0";
    tmp(32613) := x"07e0";
    tmp(32614) := x"07e0";
    tmp(32615) := x"07e0";
    tmp(32616) := x"07e0";
    tmp(32617) := x"07e0";
    tmp(32618) := x"07e0";
    tmp(32619) := x"07e0";
    tmp(32620) := x"07e0";
    tmp(32621) := x"07e0";
    tmp(32622) := x"07e0";
    tmp(32623) := x"07e0";
    tmp(32624) := x"07e0";
    tmp(32625) := x"07e0";
    tmp(32626) := x"07e0";
    tmp(32627) := x"07e0";
    tmp(32628) := x"07e0";
    tmp(32629) := x"07e0";
    tmp(32630) := x"07e0";
    tmp(32631) := x"07e0";
    tmp(32632) := x"07e0";
    tmp(32633) := x"07e0";
    tmp(32634) := x"07e0";
    tmp(32635) := x"07e0";
    tmp(32636) := x"07e0";
    tmp(32637) := x"0840";
    tmp(32638) := x"0840";
    tmp(32639) := x"0840";
    tmp(32640) := x"0000";
    tmp(32641) := x"0083";
    tmp(32642) := x"0083";
    tmp(32643) := x"0083";
    tmp(32644) := x"00a3";
    tmp(32645) := x"00a3";
    tmp(32646) := x"00a3";
    tmp(32647) := x"00a3";
    tmp(32648) := x"0083";
    tmp(32649) := x"00a3";
    tmp(32650) := x"00a4";
    tmp(32651) := x"00c4";
    tmp(32652) := x"00c4";
    tmp(32653) := x"00c5";
    tmp(32654) := x"00e5";
    tmp(32655) := x"00e5";
    tmp(32656) := x"00e5";
    tmp(32657) := x"00c5";
    tmp(32658) := x"00a4";
    tmp(32659) := x"00c4";
    tmp(32660) := x"00c4";
    tmp(32661) := x"00a3";
    tmp(32662) := x"0083";
    tmp(32663) := x"00a4";
    tmp(32664) := x"00c4";
    tmp(32665) := x"00e4";
    tmp(32666) := x"00e4";
    tmp(32667) := x"00c4";
    tmp(32668) := x"00e4";
    tmp(32669) := x"00c4";
    tmp(32670) := x"08e5";
    tmp(32671) := x"08e5";
    tmp(32672) := x"0906";
    tmp(32673) := x"0925";
    tmp(32674) := x"0925";
    tmp(32675) := x"0905";
    tmp(32676) := x"0905";
    tmp(32677) := x"0905";
    tmp(32678) := x"0905";
    tmp(32679) := x"0905";
    tmp(32680) := x"0905";
    tmp(32681) := x"0925";
    tmp(32682) := x"0905";
    tmp(32683) := x"0904";
    tmp(32684) := x"08e4";
    tmp(32685) := x"08e4";
    tmp(32686) := x"08a3";
    tmp(32687) := x"0904";
    tmp(32688) := x"0926";
    tmp(32689) := x"0946";
    tmp(32690) := x"0925";
    tmp(32691) := x"0904";
    tmp(32692) := x"1104";
    tmp(32693) := x"08c2";
    tmp(32694) := x"08c1";
    tmp(32695) := x"1121";
    tmp(32696) := x"1141";
    tmp(32697) := x"1141";
    tmp(32698) := x"1141";
    tmp(32699) := x"1140";
    tmp(32700) := x"1140";
    tmp(32701) := x"1140";
    tmp(32702) := x"1120";
    tmp(32703) := x"1120";
    tmp(32704) := x"1120";
    tmp(32705) := x"1120";
    tmp(32706) := x"1120";
    tmp(32707) := x"1120";
    tmp(32708) := x"0920";
    tmp(32709) := x"0920";
    tmp(32710) := x"0900";
    tmp(32711) := x"0900";
    tmp(32712) := x"0900";
    tmp(32713) := x"0900";
    tmp(32714) := x"0901";
    tmp(32715) := x"1101";
    tmp(32716) := x"1101";
    tmp(32717) := x"1121";
    tmp(32718) := x"1942";
    tmp(32719) := x"1942";
    tmp(32720) := x"2163";
    tmp(32721) := x"2163";
    tmp(32722) := x"2984";
    tmp(32723) := x"31a5";
    tmp(32724) := x"31c5";
    tmp(32725) := x"39e6";
    tmp(32726) := x"39e6";
    tmp(32727) := x"39e7";
    tmp(32728) := x"4207";
    tmp(32729) := x"4208";
    tmp(32730) := x"4208";
    tmp(32731) := x"4208";
    tmp(32732) := x"4208";
    tmp(32733) := x"4227";
    tmp(32734) := x"3a06";
    tmp(32735) := x"39c6";
    tmp(32736) := x"31c5";
    tmp(32737) := x"31a5";
    tmp(32738) := x"2985";
    tmp(32739) := x"2985";
    tmp(32740) := x"2985";
    tmp(32741) := x"29a5";
    tmp(32742) := x"29a5";
    tmp(32743) := x"29a5";
    tmp(32744) := x"29c5";
    tmp(32745) := x"29e5";
    tmp(32746) := x"29e5";
    tmp(32747) := x"1983";
    tmp(32748) := x"1983";
    tmp(32749) := x"1983";
    tmp(32750) := x"21a2";
    tmp(32751) := x"19a2";
    tmp(32752) := x"1981";
    tmp(32753) := x"1121";
    tmp(32754) := x"1101";
    tmp(32755) := x"1121";
    tmp(32756) := x"1121";
    tmp(32757) := x"1121";
    tmp(32758) := x"1120";
    tmp(32759) := x"1100";
    tmp(32760) := x"1100";
    tmp(32761) := x"1100";
    tmp(32762) := x"1100";
    tmp(32763) := x"1120";
    tmp(32764) := x"1120";
    tmp(32765) := x"1120";
    tmp(32766) := x"1100";
    tmp(32767) := x"1100";
    tmp(32768) := x"0900";
    tmp(32769) := x"1120";
    tmp(32770) := x"1120";
    tmp(32771) := x"1120";
    tmp(32772) := x"1140";
    tmp(32773) := x"1140";
    tmp(32774) := x"1140";
    tmp(32775) := x"1120";
    tmp(32776) := x"1121";
    tmp(32777) := x"1120";
    tmp(32778) := x"1120";
    tmp(32779) := x"1120";
    tmp(32780) := x"1920";
    tmp(32781) := x"1920";
    tmp(32782) := x"1921";
    tmp(32783) := x"1921";
    tmp(32784) := x"1921";
    tmp(32785) := x"2141";
    tmp(32786) := x"2141";
    tmp(32787) := x"2121";
    tmp(32788) := x"2121";
    tmp(32789) := x"2121";
    tmp(32790) := x"2121";
    tmp(32791) := x"2121";
    tmp(32792) := x"2121";
    tmp(32793) := x"18e1";
    tmp(32794) := x"18c1";
    tmp(32795) := x"18c1";
    tmp(32796) := x"18c1";
    tmp(32797) := x"18e1";
    tmp(32798) := x"2101";
    tmp(32799) := x"2122";
    tmp(32800) := x"2142";
    tmp(32801) := x"2142";
    tmp(32802) := x"2942";
    tmp(32803) := x"2122";
    tmp(32804) := x"2122";
    tmp(32805) := x"2122";
    tmp(32806) := x"2122";
    tmp(32807) := x"2102";
    tmp(32808) := x"2102";
    tmp(32809) := x"2102";
    tmp(32810) := x"2102";
    tmp(32811) := x"2102";
    tmp(32812) := x"20e2";
    tmp(32813) := x"20c2";
    tmp(32814) := x"20c2";
    tmp(32815) := x"20c2";
    tmp(32816) := x"20c2";
    tmp(32817) := x"18c2";
    tmp(32818) := x"20a2";
    tmp(32819) := x"20a2";
    tmp(32820) := x"18a1";
    tmp(32821) := x"18a1";
    tmp(32822) := x"18a1";
    tmp(32823) := x"18a1";
    tmp(32824) := x"18a1";
    tmp(32825) := x"1881";
    tmp(32826) := x"1881";
    tmp(32827) := x"1881";
    tmp(32828) := x"1881";
    tmp(32829) := x"1881";
    tmp(32830) := x"1881";
    tmp(32831) := x"1881";
    tmp(32832) := x"18a1";
    tmp(32833) := x"18a1";
    tmp(32834) := x"18a2";
    tmp(32835) := x"20c2";
    tmp(32836) := x"20c2";
    tmp(32837) := x"07e0";
    tmp(32838) := x"07e0";
    tmp(32839) := x"07e0";
    tmp(32840) := x"07e0";
    tmp(32841) := x"07e0";
    tmp(32842) := x"07e0";
    tmp(32843) := x"07e0";
    tmp(32844) := x"07e0";
    tmp(32845) := x"07e0";
    tmp(32846) := x"07e0";
    tmp(32847) := x"07e0";
    tmp(32848) := x"07e0";
    tmp(32849) := x"07e0";
    tmp(32850) := x"07e0";
    tmp(32851) := x"07e0";
    tmp(32852) := x"07e0";
    tmp(32853) := x"07e0";
    tmp(32854) := x"07e0";
    tmp(32855) := x"07e0";
    tmp(32856) := x"07e0";
    tmp(32857) := x"07e0";
    tmp(32858) := x"07e0";
    tmp(32859) := x"07e0";
    tmp(32860) := x"07e0";
    tmp(32861) := x"07e0";
    tmp(32862) := x"07e0";
    tmp(32863) := x"07e0";
    tmp(32864) := x"07e0";
    tmp(32865) := x"07e0";
    tmp(32866) := x"07e0";
    tmp(32867) := x"07e0";
    tmp(32868) := x"07e0";
    tmp(32869) := x"07e0";
    tmp(32870) := x"07e0";
    tmp(32871) := x"07e0";
    tmp(32872) := x"07e0";
    tmp(32873) := x"07e0";
    tmp(32874) := x"07e0";
    tmp(32875) := x"07e0";
    tmp(32876) := x"07e0";
    tmp(32877) := x"0840";
    tmp(32878) := x"0840";
    tmp(32879) := x"0840";
    tmp(32880) := x"0000";
    tmp(32881) := x"00a3";
    tmp(32882) := x"00a3";
    tmp(32883) := x"00a3";
    tmp(32884) := x"0083";
    tmp(32885) := x"0082";
    tmp(32886) := x"0062";
    tmp(32887) := x"0062";
    tmp(32888) := x"0062";
    tmp(32889) := x"0062";
    tmp(32890) := x"0062";
    tmp(32891) := x"0062";
    tmp(32892) := x"0062";
    tmp(32893) := x"0062";
    tmp(32894) := x"0062";
    tmp(32895) := x"0062";
    tmp(32896) := x"0082";
    tmp(32897) := x"00a3";
    tmp(32898) := x"00c4";
    tmp(32899) := x"00a4";
    tmp(32900) := x"00a3";
    tmp(32901) := x"00a3";
    tmp(32902) := x"0082";
    tmp(32903) := x"00a3";
    tmp(32904) := x"00c4";
    tmp(32905) := x"00c4";
    tmp(32906) := x"00c4";
    tmp(32907) := x"00c4";
    tmp(32908) := x"00e4";
    tmp(32909) := x"00c3";
    tmp(32910) := x"08e5";
    tmp(32911) := x"0905";
    tmp(32912) := x"0905";
    tmp(32913) := x"0905";
    tmp(32914) := x"0905";
    tmp(32915) := x"0905";
    tmp(32916) := x"0905";
    tmp(32917) := x"0925";
    tmp(32918) := x"0925";
    tmp(32919) := x"0905";
    tmp(32920) := x"0905";
    tmp(32921) := x"0905";
    tmp(32922) := x"08e4";
    tmp(32923) := x"08c3";
    tmp(32924) := x"08a3";
    tmp(32925) := x"08a2";
    tmp(32926) := x"0882";
    tmp(32927) := x"08e4";
    tmp(32928) := x"1187";
    tmp(32929) := x"11a7";
    tmp(32930) := x"1186";
    tmp(32931) := x"1165";
    tmp(32932) := x"1165";
    tmp(32933) := x"1122";
    tmp(32934) := x"1141";
    tmp(32935) := x"1141";
    tmp(32936) := x"1161";
    tmp(32937) := x"1141";
    tmp(32938) := x"1161";
    tmp(32939) := x"1140";
    tmp(32940) := x"1120";
    tmp(32941) := x"1120";
    tmp(32942) := x"1140";
    tmp(32943) := x"1120";
    tmp(32944) := x"1120";
    tmp(32945) := x"1120";
    tmp(32946) := x"1120";
    tmp(32947) := x"1120";
    tmp(32948) := x"0920";
    tmp(32949) := x"0920";
    tmp(32950) := x"0900";
    tmp(32951) := x"0900";
    tmp(32952) := x"0900";
    tmp(32953) := x"0900";
    tmp(32954) := x"0900";
    tmp(32955) := x"0901";
    tmp(32956) := x"1101";
    tmp(32957) := x"1121";
    tmp(32958) := x"1121";
    tmp(32959) := x"1922";
    tmp(32960) := x"1942";
    tmp(32961) := x"2143";
    tmp(32962) := x"2163";
    tmp(32963) := x"2984";
    tmp(32964) := x"31a5";
    tmp(32965) := x"31a5";
    tmp(32966) := x"31a5";
    tmp(32967) := x"39c6";
    tmp(32968) := x"39c6";
    tmp(32969) := x"39c7";
    tmp(32970) := x"39e7";
    tmp(32971) := x"39e6";
    tmp(32972) := x"39e7";
    tmp(32973) := x"39e6";
    tmp(32974) := x"31c5";
    tmp(32975) := x"31a5";
    tmp(32976) := x"3185";
    tmp(32977) := x"2984";
    tmp(32978) := x"2984";
    tmp(32979) := x"2985";
    tmp(32980) := x"2985";
    tmp(32981) := x"29a5";
    tmp(32982) := x"29c5";
    tmp(32983) := x"29c5";
    tmp(32984) := x"29e5";
    tmp(32985) := x"29c4";
    tmp(32986) := x"21a4";
    tmp(32987) := x"1963";
    tmp(32988) := x"1982";
    tmp(32989) := x"21a2";
    tmp(32990) := x"1982";
    tmp(32991) := x"1961";
    tmp(32992) := x"1141";
    tmp(32993) := x"1101";
    tmp(32994) := x"0901";
    tmp(32995) := x"1101";
    tmp(32996) := x"0901";
    tmp(32997) := x"1100";
    tmp(32998) := x"1120";
    tmp(32999) := x"1100";
    tmp(33000) := x"1100";
    tmp(33001) := x"1100";
    tmp(33002) := x"1120";
    tmp(33003) := x"1120";
    tmp(33004) := x"1120";
    tmp(33005) := x"1120";
    tmp(33006) := x"1100";
    tmp(33007) := x"1100";
    tmp(33008) := x"0900";
    tmp(33009) := x"0900";
    tmp(33010) := x"0900";
    tmp(33011) := x"1120";
    tmp(33012) := x"1120";
    tmp(33013) := x"1140";
    tmp(33014) := x"1120";
    tmp(33015) := x"1120";
    tmp(33016) := x"1120";
    tmp(33017) := x"1120";
    tmp(33018) := x"1120";
    tmp(33019) := x"1100";
    tmp(33020) := x"1100";
    tmp(33021) := x"1920";
    tmp(33022) := x"1920";
    tmp(33023) := x"1920";
    tmp(33024) := x"1921";
    tmp(33025) := x"1921";
    tmp(33026) := x"2121";
    tmp(33027) := x"2121";
    tmp(33028) := x"2121";
    tmp(33029) := x"2121";
    tmp(33030) := x"2121";
    tmp(33031) := x"2121";
    tmp(33032) := x"2121";
    tmp(33033) := x"1901";
    tmp(33034) := x"18c1";
    tmp(33035) := x"10c1";
    tmp(33036) := x"18c1";
    tmp(33037) := x"18e1";
    tmp(33038) := x"18e1";
    tmp(33039) := x"2102";
    tmp(33040) := x"2122";
    tmp(33041) := x"2122";
    tmp(33042) := x"2122";
    tmp(33043) := x"2122";
    tmp(33044) := x"2102";
    tmp(33045) := x"2102";
    tmp(33046) := x"1902";
    tmp(33047) := x"1902";
    tmp(33048) := x"1902";
    tmp(33049) := x"2102";
    tmp(33050) := x"20e2";
    tmp(33051) := x"18c2";
    tmp(33052) := x"18c2";
    tmp(33053) := x"18c2";
    tmp(33054) := x"18a2";
    tmp(33055) := x"18a1";
    tmp(33056) := x"18a1";
    tmp(33057) := x"18a1";
    tmp(33058) := x"18a1";
    tmp(33059) := x"18a1";
    tmp(33060) := x"1881";
    tmp(33061) := x"1881";
    tmp(33062) := x"1881";
    tmp(33063) := x"1881";
    tmp(33064) := x"1881";
    tmp(33065) := x"1881";
    tmp(33066) := x"1881";
    tmp(33067) := x"1881";
    tmp(33068) := x"1881";
    tmp(33069) := x"1881";
    tmp(33070) := x"1881";
    tmp(33071) := x"1881";
    tmp(33072) := x"1881";
    tmp(33073) := x"1881";
    tmp(33074) := x"1881";
    tmp(33075) := x"18a1";
    tmp(33076) := x"18a1";
    tmp(33077) := x"07e0";
    tmp(33078) := x"07e0";
    tmp(33079) := x"07e0";
    tmp(33080) := x"07e0";
    tmp(33081) := x"07e0";
    tmp(33082) := x"07e0";
    tmp(33083) := x"07e0";
    tmp(33084) := x"07e0";
    tmp(33085) := x"07e0";
    tmp(33086) := x"07e0";
    tmp(33087) := x"07e0";
    tmp(33088) := x"07e0";
    tmp(33089) := x"07e0";
    tmp(33090) := x"07e0";
    tmp(33091) := x"07e0";
    tmp(33092) := x"07e0";
    tmp(33093) := x"07e0";
    tmp(33094) := x"07e0";
    tmp(33095) := x"07e0";
    tmp(33096) := x"07e0";
    tmp(33097) := x"07e0";
    tmp(33098) := x"07e0";
    tmp(33099) := x"07e0";
    tmp(33100) := x"07e0";
    tmp(33101) := x"07e0";
    tmp(33102) := x"07e0";
    tmp(33103) := x"07e0";
    tmp(33104) := x"07e0";
    tmp(33105) := x"07e0";
    tmp(33106) := x"07e0";
    tmp(33107) := x"07e0";
    tmp(33108) := x"07e0";
    tmp(33109) := x"07e0";
    tmp(33110) := x"07e0";
    tmp(33111) := x"07e0";
    tmp(33112) := x"07e0";
    tmp(33113) := x"07e0";
    tmp(33114) := x"07e0";
    tmp(33115) := x"07e0";
    tmp(33116) := x"07e0";
    tmp(33117) := x"0840";
    tmp(33118) := x"0840";
    tmp(33119) := x"0840";
    tmp(33120) := x"0000";
    tmp(33121) := x"0083";
    tmp(33122) := x"0083";
    tmp(33123) := x"0082";
    tmp(33124) := x"0082";
    tmp(33125) := x"0082";
    tmp(33126) := x"0083";
    tmp(33127) := x"0083";
    tmp(33128) := x"0083";
    tmp(33129) := x"0083";
    tmp(33130) := x"0062";
    tmp(33131) := x"0062";
    tmp(33132) := x"0062";
    tmp(33133) := x"0062";
    tmp(33134) := x"0062";
    tmp(33135) := x"0062";
    tmp(33136) := x"0082";
    tmp(33137) := x"00a3";
    tmp(33138) := x"00c4";
    tmp(33139) := x"00c4";
    tmp(33140) := x"00c4";
    tmp(33141) := x"08e4";
    tmp(33142) := x"00c4";
    tmp(33143) := x"00a3";
    tmp(33144) := x"00c4";
    tmp(33145) := x"0905";
    tmp(33146) := x"0906";
    tmp(33147) := x"0905";
    tmp(33148) := x"08e5";
    tmp(33149) := x"00c4";
    tmp(33150) := x"08e5";
    tmp(33151) := x"0905";
    tmp(33152) := x"0905";
    tmp(33153) := x"0905";
    tmp(33154) := x"08e5";
    tmp(33155) := x"08e4";
    tmp(33156) := x"0905";
    tmp(33157) := x"0905";
    tmp(33158) := x"0905";
    tmp(33159) := x"0905";
    tmp(33160) := x"0904";
    tmp(33161) := x"0904";
    tmp(33162) := x"08e4";
    tmp(33163) := x"08c3";
    tmp(33164) := x"08a2";
    tmp(33165) := x"08a2";
    tmp(33166) := x"08a3";
    tmp(33167) := x"11a7";
    tmp(33168) := x"11a8";
    tmp(33169) := x"1186";
    tmp(33170) := x"1165";
    tmp(33171) := x"1185";
    tmp(33172) := x"11a4";
    tmp(33173) := x"1141";
    tmp(33174) := x"1141";
    tmp(33175) := x"1141";
    tmp(33176) := x"1141";
    tmp(33177) := x"1141";
    tmp(33178) := x"1140";
    tmp(33179) := x"1141";
    tmp(33180) := x"1140";
    tmp(33181) := x"1140";
    tmp(33182) := x"1140";
    tmp(33183) := x"1140";
    tmp(33184) := x"1140";
    tmp(33185) := x"1140";
    tmp(33186) := x"1120";
    tmp(33187) := x"1120";
    tmp(33188) := x"1120";
    tmp(33189) := x"0920";
    tmp(33190) := x"0920";
    tmp(33191) := x"0900";
    tmp(33192) := x"0900";
    tmp(33193) := x"0900";
    tmp(33194) := x"0900";
    tmp(33195) := x"08e1";
    tmp(33196) := x"1101";
    tmp(33197) := x"1101";
    tmp(33198) := x"1101";
    tmp(33199) := x"1101";
    tmp(33200) := x"1922";
    tmp(33201) := x"1942";
    tmp(33202) := x"2163";
    tmp(33203) := x"2163";
    tmp(33204) := x"2984";
    tmp(33205) := x"2984";
    tmp(33206) := x"2984";
    tmp(33207) := x"3185";
    tmp(33208) := x"3185";
    tmp(33209) := x"31a6";
    tmp(33210) := x"39c6";
    tmp(33211) := x"31a6";
    tmp(33212) := x"39a5";
    tmp(33213) := x"31a5";
    tmp(33214) := x"2984";
    tmp(33215) := x"2964";
    tmp(33216) := x"2964";
    tmp(33217) := x"2964";
    tmp(33218) := x"2984";
    tmp(33219) := x"2985";
    tmp(33220) := x"29a5";
    tmp(33221) := x"31c5";
    tmp(33222) := x"29c5";
    tmp(33223) := x"29c5";
    tmp(33224) := x"29c4";
    tmp(33225) := x"21a4";
    tmp(33226) := x"1963";
    tmp(33227) := x"1942";
    tmp(33228) := x"1982";
    tmp(33229) := x"1982";
    tmp(33230) := x"1961";
    tmp(33231) := x"1141";
    tmp(33232) := x"1121";
    tmp(33233) := x"0900";
    tmp(33234) := x"0901";
    tmp(33235) := x"1101";
    tmp(33236) := x"1101";
    tmp(33237) := x"1100";
    tmp(33238) := x"1100";
    tmp(33239) := x"1100";
    tmp(33240) := x"0900";
    tmp(33241) := x"1100";
    tmp(33242) := x"1120";
    tmp(33243) := x"1120";
    tmp(33244) := x"1120";
    tmp(33245) := x"1120";
    tmp(33246) := x"1120";
    tmp(33247) := x"1120";
    tmp(33248) := x"0900";
    tmp(33249) := x"0900";
    tmp(33250) := x"0900";
    tmp(33251) := x"1120";
    tmp(33252) := x"1120";
    tmp(33253) := x"1120";
    tmp(33254) := x"1120";
    tmp(33255) := x"1120";
    tmp(33256) := x"1120";
    tmp(33257) := x"1120";
    tmp(33258) := x"1120";
    tmp(33259) := x"1100";
    tmp(33260) := x"1100";
    tmp(33261) := x"1100";
    tmp(33262) := x"1920";
    tmp(33263) := x"1900";
    tmp(33264) := x"1901";
    tmp(33265) := x"1921";
    tmp(33266) := x"1921";
    tmp(33267) := x"1921";
    tmp(33268) := x"2121";
    tmp(33269) := x"2121";
    tmp(33270) := x"2121";
    tmp(33271) := x"1901";
    tmp(33272) := x"1901";
    tmp(33273) := x"1901";
    tmp(33274) := x"18c1";
    tmp(33275) := x"10c1";
    tmp(33276) := x"10a1";
    tmp(33277) := x"10c1";
    tmp(33278) := x"18c1";
    tmp(33279) := x"18e1";
    tmp(33280) := x"2102";
    tmp(33281) := x"2102";
    tmp(33282) := x"18e1";
    tmp(33283) := x"18e1";
    tmp(33284) := x"18e1";
    tmp(33285) := x"18e1";
    tmp(33286) := x"18c1";
    tmp(33287) := x"18e1";
    tmp(33288) := x"18c1";
    tmp(33289) := x"18c1";
    tmp(33290) := x"18c1";
    tmp(33291) := x"18c1";
    tmp(33292) := x"18a1";
    tmp(33293) := x"18a1";
    tmp(33294) := x"18a1";
    tmp(33295) := x"18a1";
    tmp(33296) := x"1881";
    tmp(33297) := x"1881";
    tmp(33298) := x"1881";
    tmp(33299) := x"1881";
    tmp(33300) := x"1881";
    tmp(33301) := x"1881";
    tmp(33302) := x"1881";
    tmp(33303) := x"1881";
    tmp(33304) := x"1881";
    tmp(33305) := x"1861";
    tmp(33306) := x"1061";
    tmp(33307) := x"1061";
    tmp(33308) := x"1061";
    tmp(33309) := x"1061";
    tmp(33310) := x"1061";
    tmp(33311) := x"1061";
    tmp(33312) := x"1061";
    tmp(33313) := x"1081";
    tmp(33314) := x"1081";
    tmp(33315) := x"1081";
    tmp(33316) := x"1881";
    tmp(33317) := x"07e0";
    tmp(33318) := x"07e0";
    tmp(33319) := x"07e0";
    tmp(33320) := x"07e0";
    tmp(33321) := x"07e0";
    tmp(33322) := x"07e0";
    tmp(33323) := x"07e0";
    tmp(33324) := x"07e0";
    tmp(33325) := x"07e0";
    tmp(33326) := x"07e0";
    tmp(33327) := x"07e0";
    tmp(33328) := x"07e0";
    tmp(33329) := x"07e0";
    tmp(33330) := x"07e0";
    tmp(33331) := x"07e0";
    tmp(33332) := x"07e0";
    tmp(33333) := x"07e0";
    tmp(33334) := x"07e0";
    tmp(33335) := x"07e0";
    tmp(33336) := x"07e0";
    tmp(33337) := x"07e0";
    tmp(33338) := x"07e0";
    tmp(33339) := x"07e0";
    tmp(33340) := x"07e0";
    tmp(33341) := x"07e0";
    tmp(33342) := x"07e0";
    tmp(33343) := x"07e0";
    tmp(33344) := x"07e0";
    tmp(33345) := x"07e0";
    tmp(33346) := x"07e0";
    tmp(33347) := x"07e0";
    tmp(33348) := x"07e0";
    tmp(33349) := x"07e0";
    tmp(33350) := x"07e0";
    tmp(33351) := x"07e0";
    tmp(33352) := x"07e0";
    tmp(33353) := x"07e0";
    tmp(33354) := x"07e0";
    tmp(33355) := x"07e0";
    tmp(33356) := x"07e0";
    tmp(33357) := x"0840";
    tmp(33358) := x"0840";
    tmp(33359) := x"0840";
    tmp(33360) := x"0000";
    tmp(33361) := x"0082";
    tmp(33362) := x"0082";
    tmp(33363) := x"0082";
    tmp(33364) := x"0062";
    tmp(33365) := x"0062";
    tmp(33366) := x"0062";
    tmp(33367) := x"0062";
    tmp(33368) := x"0062";
    tmp(33369) := x"0083";
    tmp(33370) := x"0083";
    tmp(33371) := x"00a3";
    tmp(33372) := x"00c4";
    tmp(33373) := x"00c4";
    tmp(33374) := x"00c4";
    tmp(33375) := x"00c4";
    tmp(33376) := x"00c4";
    tmp(33377) := x"00c3";
    tmp(33378) := x"00c4";
    tmp(33379) := x"00e5";
    tmp(33380) := x"00e5";
    tmp(33381) := x"00e5";
    tmp(33382) := x"00e4";
    tmp(33383) := x"00c4";
    tmp(33384) := x"00a3";
    tmp(33385) := x"00c4";
    tmp(33386) := x"00c4";
    tmp(33387) := x"00e5";
    tmp(33388) := x"0926";
    tmp(33389) := x"0905";
    tmp(33390) := x"0906";
    tmp(33391) := x"0926";
    tmp(33392) := x"0906";
    tmp(33393) := x"0906";
    tmp(33394) := x"0905";
    tmp(33395) := x"0925";
    tmp(33396) := x"0925";
    tmp(33397) := x"0925";
    tmp(33398) := x"0925";
    tmp(33399) := x"0925";
    tmp(33400) := x"0945";
    tmp(33401) := x"0925";
    tmp(33402) := x"0925";
    tmp(33403) := x"0904";
    tmp(33404) := x"08e4";
    tmp(33405) := x"0904";
    tmp(33406) := x"0925";
    tmp(33407) := x"11c8";
    tmp(33408) := x"1186";
    tmp(33409) := x"1145";
    tmp(33410) := x"1124";
    tmp(33411) := x"11a4";
    tmp(33412) := x"1161";
    tmp(33413) := x"1141";
    tmp(33414) := x"1141";
    tmp(33415) := x"1141";
    tmp(33416) := x"1141";
    tmp(33417) := x"1141";
    tmp(33418) := x"1141";
    tmp(33419) := x"1161";
    tmp(33420) := x"1140";
    tmp(33421) := x"1141";
    tmp(33422) := x"1140";
    tmp(33423) := x"1140";
    tmp(33424) := x"1140";
    tmp(33425) := x"1140";
    tmp(33426) := x"1140";
    tmp(33427) := x"1120";
    tmp(33428) := x"1120";
    tmp(33429) := x"0920";
    tmp(33430) := x"0920";
    tmp(33431) := x"0920";
    tmp(33432) := x"0900";
    tmp(33433) := x"0900";
    tmp(33434) := x"0900";
    tmp(33435) := x"0901";
    tmp(33436) := x"0901";
    tmp(33437) := x"1101";
    tmp(33438) := x"1101";
    tmp(33439) := x"1101";
    tmp(33440) := x"1122";
    tmp(33441) := x"1922";
    tmp(33442) := x"1942";
    tmp(33443) := x"2143";
    tmp(33444) := x"2143";
    tmp(33445) := x"2163";
    tmp(33446) := x"2943";
    tmp(33447) := x"2964";
    tmp(33448) := x"2964";
    tmp(33449) := x"3185";
    tmp(33450) := x"3185";
    tmp(33451) := x"3185";
    tmp(33452) := x"2964";
    tmp(33453) := x"2964";
    tmp(33454) := x"2943";
    tmp(33455) := x"2943";
    tmp(33456) := x"2944";
    tmp(33457) := x"2964";
    tmp(33458) := x"2985";
    tmp(33459) := x"31a5";
    tmp(33460) := x"31c5";
    tmp(33461) := x"29a5";
    tmp(33462) := x"29a4";
    tmp(33463) := x"29a4";
    tmp(33464) := x"21a3";
    tmp(33465) := x"2183";
    tmp(33466) := x"1942";
    tmp(33467) := x"1962";
    tmp(33468) := x"1962";
    tmp(33469) := x"1961";
    tmp(33470) := x"1141";
    tmp(33471) := x"1141";
    tmp(33472) := x"1121";
    tmp(33473) := x"0900";
    tmp(33474) := x"0901";
    tmp(33475) := x"1101";
    tmp(33476) := x"1100";
    tmp(33477) := x"0900";
    tmp(33478) := x"1100";
    tmp(33479) := x"1100";
    tmp(33480) := x"1100";
    tmp(33481) := x"1100";
    tmp(33482) := x"1100";
    tmp(33483) := x"1120";
    tmp(33484) := x"1121";
    tmp(33485) := x"1121";
    tmp(33486) := x"1120";
    tmp(33487) := x"1120";
    tmp(33488) := x"0900";
    tmp(33489) := x"0900";
    tmp(33490) := x"0900";
    tmp(33491) := x"0900";
    tmp(33492) := x"1120";
    tmp(33493) := x"1120";
    tmp(33494) := x"1120";
    tmp(33495) := x"1120";
    tmp(33496) := x"1100";
    tmp(33497) := x"1100";
    tmp(33498) := x"1100";
    tmp(33499) := x"1100";
    tmp(33500) := x"1120";
    tmp(33501) := x"1100";
    tmp(33502) := x"1100";
    tmp(33503) := x"1900";
    tmp(33504) := x"1900";
    tmp(33505) := x"1901";
    tmp(33506) := x"1901";
    tmp(33507) := x"1901";
    tmp(33508) := x"1901";
    tmp(33509) := x"2101";
    tmp(33510) := x"1901";
    tmp(33511) := x"1901";
    tmp(33512) := x"1901";
    tmp(33513) := x"18e1";
    tmp(33514) := x"18c1";
    tmp(33515) := x"10a1";
    tmp(33516) := x"10a1";
    tmp(33517) := x"10a1";
    tmp(33518) := x"10a1";
    tmp(33519) := x"18c1";
    tmp(33520) := x"18c1";
    tmp(33521) := x"18c1";
    tmp(33522) := x"18c1";
    tmp(33523) := x"18c1";
    tmp(33524) := x"18c1";
    tmp(33525) := x"18a1";
    tmp(33526) := x"18a1";
    tmp(33527) := x"18a1";
    tmp(33528) := x"18a1";
    tmp(33529) := x"18a1";
    tmp(33530) := x"18a1";
    tmp(33531) := x"18a1";
    tmp(33532) := x"18a1";
    tmp(33533) := x"1081";
    tmp(33534) := x"1081";
    tmp(33535) := x"1081";
    tmp(33536) := x"1081";
    tmp(33537) := x"1081";
    tmp(33538) := x"1881";
    tmp(33539) := x"1881";
    tmp(33540) := x"1081";
    tmp(33541) := x"1061";
    tmp(33542) := x"1061";
    tmp(33543) := x"1061";
    tmp(33544) := x"1061";
    tmp(33545) := x"1061";
    tmp(33546) := x"1061";
    tmp(33547) := x"1061";
    tmp(33548) := x"1061";
    tmp(33549) := x"1061";
    tmp(33550) := x"1061";
    tmp(33551) := x"1061";
    tmp(33552) := x"1061";
    tmp(33553) := x"1061";
    tmp(33554) := x"1061";
    tmp(33555) := x"1061";
    tmp(33556) := x"1061";
    tmp(33557) := x"07e0";
    tmp(33558) := x"07e0";
    tmp(33559) := x"07e0";
    tmp(33560) := x"07e0";
    tmp(33561) := x"07e0";
    tmp(33562) := x"07e0";
    tmp(33563) := x"07e0";
    tmp(33564) := x"07e0";
    tmp(33565) := x"07e0";
    tmp(33566) := x"07e0";
    tmp(33567) := x"07e0";
    tmp(33568) := x"07e0";
    tmp(33569) := x"07e0";
    tmp(33570) := x"07e0";
    tmp(33571) := x"07e0";
    tmp(33572) := x"07e0";
    tmp(33573) := x"07e0";
    tmp(33574) := x"07e0";
    tmp(33575) := x"07e0";
    tmp(33576) := x"07e0";
    tmp(33577) := x"07e0";
    tmp(33578) := x"07e0";
    tmp(33579) := x"07e0";
    tmp(33580) := x"07e0";
    tmp(33581) := x"07e0";
    tmp(33582) := x"07e0";
    tmp(33583) := x"07e0";
    tmp(33584) := x"07e0";
    tmp(33585) := x"07e0";
    tmp(33586) := x"07e0";
    tmp(33587) := x"07e0";
    tmp(33588) := x"07e0";
    tmp(33589) := x"07e0";
    tmp(33590) := x"07e0";
    tmp(33591) := x"07e0";
    tmp(33592) := x"07e0";
    tmp(33593) := x"07e0";
    tmp(33594) := x"07e0";
    tmp(33595) := x"07e0";
    tmp(33596) := x"07e0";
    tmp(33597) := x"0840";
    tmp(33598) := x"0840";
    tmp(33599) := x"0840";
    tmp(33600) := x"0000";
    tmp(33601) := x"0083";
    tmp(33602) := x"0082";
    tmp(33603) := x"0082";
    tmp(33604) := x"0082";
    tmp(33605) := x"0062";
    tmp(33606) := x"0083";
    tmp(33607) := x"00a4";
    tmp(33608) := x"00c4";
    tmp(33609) := x"00e5";
    tmp(33610) := x"00e5";
    tmp(33611) := x"00e5";
    tmp(33612) := x"00e5";
    tmp(33613) := x"00e5";
    tmp(33614) := x"00c4";
    tmp(33615) := x"00c4";
    tmp(33616) := x"00e4";
    tmp(33617) := x"00e5";
    tmp(33618) := x"0105";
    tmp(33619) := x"0105";
    tmp(33620) := x"0105";
    tmp(33621) := x"00e5";
    tmp(33622) := x"00e4";
    tmp(33623) := x"00c4";
    tmp(33624) := x"00a3";
    tmp(33625) := x"00a3";
    tmp(33626) := x"00c4";
    tmp(33627) := x"08e5";
    tmp(33628) := x"0905";
    tmp(33629) := x"08c4";
    tmp(33630) := x"08e4";
    tmp(33631) := x"0905";
    tmp(33632) := x"0947";
    tmp(33633) := x"0926";
    tmp(33634) := x"0926";
    tmp(33635) := x"0947";
    tmp(33636) := x"0967";
    tmp(33637) := x"0946";
    tmp(33638) := x"0966";
    tmp(33639) := x"0986";
    tmp(33640) := x"0987";
    tmp(33641) := x"0967";
    tmp(33642) := x"0926";
    tmp(33643) := x"0905";
    tmp(33644) := x"0946";
    tmp(33645) := x"11a7";
    tmp(33646) := x"11e9";
    tmp(33647) := x"1a8b";
    tmp(33648) := x"11e8";
    tmp(33649) := x"1185";
    tmp(33650) := x"1183";
    tmp(33651) := x"1161";
    tmp(33652) := x"1141";
    tmp(33653) := x"1140";
    tmp(33654) := x"1140";
    tmp(33655) := x"1140";
    tmp(33656) := x"1141";
    tmp(33657) := x"1140";
    tmp(33658) := x"1161";
    tmp(33659) := x"1161";
    tmp(33660) := x"1161";
    tmp(33661) := x"1141";
    tmp(33662) := x"1161";
    tmp(33663) := x"1140";
    tmp(33664) := x"1140";
    tmp(33665) := x"1140";
    tmp(33666) := x"1140";
    tmp(33667) := x"1140";
    tmp(33668) := x"1120";
    tmp(33669) := x"1120";
    tmp(33670) := x"0920";
    tmp(33671) := x"0900";
    tmp(33672) := x"0900";
    tmp(33673) := x"0900";
    tmp(33674) := x"0900";
    tmp(33675) := x"08e0";
    tmp(33676) := x"08e1";
    tmp(33677) := x"08e1";
    tmp(33678) := x"1101";
    tmp(33679) := x"1101";
    tmp(33680) := x"1101";
    tmp(33681) := x"1922";
    tmp(33682) := x"1922";
    tmp(33683) := x"1922";
    tmp(33684) := x"1923";
    tmp(33685) := x"2123";
    tmp(33686) := x"2143";
    tmp(33687) := x"2143";
    tmp(33688) := x"2944";
    tmp(33689) := x"2964";
    tmp(33690) := x"2964";
    tmp(33691) := x"2964";
    tmp(33692) := x"2143";
    tmp(33693) := x"2123";
    tmp(33694) := x"2123";
    tmp(33695) := x"2943";
    tmp(33696) := x"2964";
    tmp(33697) := x"2964";
    tmp(33698) := x"31a5";
    tmp(33699) := x"31a5";
    tmp(33700) := x"29a4";
    tmp(33701) := x"2984";
    tmp(33702) := x"2183";
    tmp(33703) := x"2183";
    tmp(33704) := x"2162";
    tmp(33705) := x"1962";
    tmp(33706) := x"1942";
    tmp(33707) := x"1961";
    tmp(33708) := x"1941";
    tmp(33709) := x"1141";
    tmp(33710) := x"1121";
    tmp(33711) := x"1121";
    tmp(33712) := x"0901";
    tmp(33713) := x"0900";
    tmp(33714) := x"0900";
    tmp(33715) := x"1100";
    tmp(33716) := x"1100";
    tmp(33717) := x"1100";
    tmp(33718) := x"1100";
    tmp(33719) := x"1100";
    tmp(33720) := x"1100";
    tmp(33721) := x"1100";
    tmp(33722) := x"1100";
    tmp(33723) := x"1100";
    tmp(33724) := x"1121";
    tmp(33725) := x"1121";
    tmp(33726) := x"1120";
    tmp(33727) := x"1120";
    tmp(33728) := x"1120";
    tmp(33729) := x"0920";
    tmp(33730) := x"0920";
    tmp(33731) := x"0900";
    tmp(33732) := x"0900";
    tmp(33733) := x"1120";
    tmp(33734) := x"1120";
    tmp(33735) := x"1120";
    tmp(33736) := x"1120";
    tmp(33737) := x"1100";
    tmp(33738) := x"1100";
    tmp(33739) := x"1100";
    tmp(33740) := x"1100";
    tmp(33741) := x"1100";
    tmp(33742) := x"1100";
    tmp(33743) := x"1100";
    tmp(33744) := x"1900";
    tmp(33745) := x"1900";
    tmp(33746) := x"1901";
    tmp(33747) := x"1901";
    tmp(33748) := x"1901";
    tmp(33749) := x"2121";
    tmp(33750) := x"1901";
    tmp(33751) := x"1901";
    tmp(33752) := x"1901";
    tmp(33753) := x"18e1";
    tmp(33754) := x"18c1";
    tmp(33755) := x"10a1";
    tmp(33756) := x"10a1";
    tmp(33757) := x"10a0";
    tmp(33758) := x"10a0";
    tmp(33759) := x"10a1";
    tmp(33760) := x"10a1";
    tmp(33761) := x"10a1";
    tmp(33762) := x"10a1";
    tmp(33763) := x"10a1";
    tmp(33764) := x"10a1";
    tmp(33765) := x"10a1";
    tmp(33766) := x"10a1";
    tmp(33767) := x"10a1";
    tmp(33768) := x"10a1";
    tmp(33769) := x"1081";
    tmp(33770) := x"1081";
    tmp(33771) := x"1081";
    tmp(33772) := x"1081";
    tmp(33773) := x"1081";
    tmp(33774) := x"1081";
    tmp(33775) := x"1081";
    tmp(33776) := x"1081";
    tmp(33777) := x"1081";
    tmp(33778) := x"1061";
    tmp(33779) := x"1061";
    tmp(33780) := x"1061";
    tmp(33781) := x"1061";
    tmp(33782) := x"1061";
    tmp(33783) := x"1061";
    tmp(33784) := x"1061";
    tmp(33785) := x"1061";
    tmp(33786) := x"1061";
    tmp(33787) := x"1061";
    tmp(33788) := x"1061";
    tmp(33789) := x"1061";
    tmp(33790) := x"1061";
    tmp(33791) := x"1061";
    tmp(33792) := x"1060";
    tmp(33793) := x"1060";
    tmp(33794) := x"1060";
    tmp(33795) := x"1060";
    tmp(33796) := x"1060";
    tmp(33797) := x"07e0";
    tmp(33798) := x"07e0";
    tmp(33799) := x"07e0";
    tmp(33800) := x"07e0";
    tmp(33801) := x"07e0";
    tmp(33802) := x"07e0";
    tmp(33803) := x"07e0";
    tmp(33804) := x"07e0";
    tmp(33805) := x"07e0";
    tmp(33806) := x"07e0";
    tmp(33807) := x"07e0";
    tmp(33808) := x"07e0";
    tmp(33809) := x"07e0";
    tmp(33810) := x"07e0";
    tmp(33811) := x"07e0";
    tmp(33812) := x"07e0";
    tmp(33813) := x"07e0";
    tmp(33814) := x"07e0";
    tmp(33815) := x"07e0";
    tmp(33816) := x"07e0";
    tmp(33817) := x"07e0";
    tmp(33818) := x"07e0";
    tmp(33819) := x"07e0";
    tmp(33820) := x"07e0";
    tmp(33821) := x"07e0";
    tmp(33822) := x"07e0";
    tmp(33823) := x"07e0";
    tmp(33824) := x"07e0";
    tmp(33825) := x"07e0";
    tmp(33826) := x"07e0";
    tmp(33827) := x"07e0";
    tmp(33828) := x"07e0";
    tmp(33829) := x"07e0";
    tmp(33830) := x"07e0";
    tmp(33831) := x"07e0";
    tmp(33832) := x"07e0";
    tmp(33833) := x"07e0";
    tmp(33834) := x"07e0";
    tmp(33835) := x"07e0";
    tmp(33836) := x"07e0";
    tmp(33837) := x"0840";
    tmp(33838) := x"0840";
    tmp(33839) := x"0840";
    tmp(33840) := x"0000";
    tmp(33841) := x"00a3";
    tmp(33842) := x"00a3";
    tmp(33843) := x"00a2";
    tmp(33844) := x"00a3";
    tmp(33845) := x"00a4";
    tmp(33846) := x"00e5";
    tmp(33847) := x"0105";
    tmp(33848) := x"0125";
    tmp(33849) := x"0105";
    tmp(33850) := x"0105";
    tmp(33851) := x"0105";
    tmp(33852) := x"00e5";
    tmp(33853) := x"00e4";
    tmp(33854) := x"00e4";
    tmp(33855) := x"0105";
    tmp(33856) := x"0105";
    tmp(33857) := x"0105";
    tmp(33858) := x"0105";
    tmp(33859) := x"0105";
    tmp(33860) := x"0105";
    tmp(33861) := x"0105";
    tmp(33862) := x"00e5";
    tmp(33863) := x"00e4";
    tmp(33864) := x"00a3";
    tmp(33865) := x"08c3";
    tmp(33866) := x"08c4";
    tmp(33867) := x"08e5";
    tmp(33868) := x"08e4";
    tmp(33869) := x"08c4";
    tmp(33870) := x"08c4";
    tmp(33871) := x"0905";
    tmp(33872) := x"08e5";
    tmp(33873) := x"0905";
    tmp(33874) := x"0926";
    tmp(33875) := x"0947";
    tmp(33876) := x"0946";
    tmp(33877) := x"0947";
    tmp(33878) := x"0987";
    tmp(33879) := x"0987";
    tmp(33880) := x"0925";
    tmp(33881) := x"08c4";
    tmp(33882) := x"08e5";
    tmp(33883) := x"0967";
    tmp(33884) := x"0987";
    tmp(33885) := x"122a";
    tmp(33886) := x"1a6b";
    tmp(33887) := x"11e8";
    tmp(33888) := x"11e7";
    tmp(33889) := x"11a3";
    tmp(33890) := x"1141";
    tmp(33891) := x"1141";
    tmp(33892) := x"1140";
    tmp(33893) := x"1140";
    tmp(33894) := x"1140";
    tmp(33895) := x"1141";
    tmp(33896) := x"1141";
    tmp(33897) := x"1161";
    tmp(33898) := x"1161";
    tmp(33899) := x"1161";
    tmp(33900) := x"1161";
    tmp(33901) := x"1161";
    tmp(33902) := x"1161";
    tmp(33903) := x"1161";
    tmp(33904) := x"1140";
    tmp(33905) := x"1120";
    tmp(33906) := x"1140";
    tmp(33907) := x"1140";
    tmp(33908) := x"1140";
    tmp(33909) := x"1120";
    tmp(33910) := x"0920";
    tmp(33911) := x"0900";
    tmp(33912) := x"0900";
    tmp(33913) := x"0900";
    tmp(33914) := x"08e0";
    tmp(33915) := x"08e0";
    tmp(33916) := x"08e0";
    tmp(33917) := x"08e1";
    tmp(33918) := x"1101";
    tmp(33919) := x"1101";
    tmp(33920) := x"1101";
    tmp(33921) := x"1101";
    tmp(33922) := x"1102";
    tmp(33923) := x"1922";
    tmp(33924) := x"1902";
    tmp(33925) := x"1902";
    tmp(33926) := x"1922";
    tmp(33927) := x"1923";
    tmp(33928) := x"2123";
    tmp(33929) := x"2143";
    tmp(33930) := x"2143";
    tmp(33931) := x"2123";
    tmp(33932) := x"2123";
    tmp(33933) := x"2123";
    tmp(33934) := x"2123";
    tmp(33935) := x"2943";
    tmp(33936) := x"2964";
    tmp(33937) := x"3184";
    tmp(33938) := x"31a4";
    tmp(33939) := x"2984";
    tmp(33940) := x"2963";
    tmp(33941) := x"2163";
    tmp(33942) := x"2162";
    tmp(33943) := x"1962";
    tmp(33944) := x"1962";
    tmp(33945) := x"1942";
    tmp(33946) := x"1941";
    tmp(33947) := x"1941";
    tmp(33948) := x"1121";
    tmp(33949) := x"1121";
    tmp(33950) := x"1121";
    tmp(33951) := x"1121";
    tmp(33952) := x"0900";
    tmp(33953) := x"0900";
    tmp(33954) := x"0900";
    tmp(33955) := x"1100";
    tmp(33956) := x"10e0";
    tmp(33957) := x"1100";
    tmp(33958) := x"1100";
    tmp(33959) := x"1100";
    tmp(33960) := x"1100";
    tmp(33961) := x"10e0";
    tmp(33962) := x"1100";
    tmp(33963) := x"1100";
    tmp(33964) := x"1120";
    tmp(33965) := x"1121";
    tmp(33966) := x"1141";
    tmp(33967) := x"1140";
    tmp(33968) := x"1120";
    tmp(33969) := x"0920";
    tmp(33970) := x"0900";
    tmp(33971) := x"0900";
    tmp(33972) := x"0900";
    tmp(33973) := x"0900";
    tmp(33974) := x"1120";
    tmp(33975) := x"1100";
    tmp(33976) := x"1120";
    tmp(33977) := x"1100";
    tmp(33978) := x"1100";
    tmp(33979) := x"10e0";
    tmp(33980) := x"1100";
    tmp(33981) := x"1100";
    tmp(33982) := x"1100";
    tmp(33983) := x"1100";
    tmp(33984) := x"1900";
    tmp(33985) := x"1900";
    tmp(33986) := x"18e0";
    tmp(33987) := x"1901";
    tmp(33988) := x"18e1";
    tmp(33989) := x"1901";
    tmp(33990) := x"1901";
    tmp(33991) := x"18e1";
    tmp(33992) := x"18e1";
    tmp(33993) := x"18c1";
    tmp(33994) := x"10c1";
    tmp(33995) := x"10a1";
    tmp(33996) := x"10a0";
    tmp(33997) := x"1080";
    tmp(33998) := x"1080";
    tmp(33999) := x"1080";
    tmp(34000) := x"1080";
    tmp(34001) := x"1080";
    tmp(34002) := x"1080";
    tmp(34003) := x"1080";
    tmp(34004) := x"1080";
    tmp(34005) := x"1080";
    tmp(34006) := x"1080";
    tmp(34007) := x"1081";
    tmp(34008) := x"1081";
    tmp(34009) := x"1081";
    tmp(34010) := x"1081";
    tmp(34011) := x"1081";
    tmp(34012) := x"1081";
    tmp(34013) := x"1061";
    tmp(34014) := x"1061";
    tmp(34015) := x"1061";
    tmp(34016) := x"1061";
    tmp(34017) := x"1061";
    tmp(34018) := x"1061";
    tmp(34019) := x"1061";
    tmp(34020) := x"1061";
    tmp(34021) := x"1061";
    tmp(34022) := x"1061";
    tmp(34023) := x"1061";
    tmp(34024) := x"1061";
    tmp(34025) := x"1061";
    tmp(34026) := x"1061";
    tmp(34027) := x"1061";
    tmp(34028) := x"1060";
    tmp(34029) := x"1060";
    tmp(34030) := x"1040";
    tmp(34031) := x"1040";
    tmp(34032) := x"1040";
    tmp(34033) := x"1040";
    tmp(34034) := x"1040";
    tmp(34035) := x"1040";
    tmp(34036) := x"1040";
    tmp(34037) := x"07e0";
    tmp(34038) := x"07e0";
    tmp(34039) := x"07e0";
    tmp(34040) := x"07e0";
    tmp(34041) := x"07e0";
    tmp(34042) := x"07e0";
    tmp(34043) := x"07e0";
    tmp(34044) := x"07e0";
    tmp(34045) := x"07e0";
    tmp(34046) := x"07e0";
    tmp(34047) := x"07e0";
    tmp(34048) := x"07e0";
    tmp(34049) := x"07e0";
    tmp(34050) := x"07e0";
    tmp(34051) := x"07e0";
    tmp(34052) := x"07e0";
    tmp(34053) := x"07e0";
    tmp(34054) := x"07e0";
    tmp(34055) := x"07e0";
    tmp(34056) := x"07e0";
    tmp(34057) := x"07e0";
    tmp(34058) := x"07e0";
    tmp(34059) := x"07e0";
    tmp(34060) := x"07e0";
    tmp(34061) := x"07e0";
    tmp(34062) := x"07e0";
    tmp(34063) := x"07e0";
    tmp(34064) := x"07e0";
    tmp(34065) := x"07e0";
    tmp(34066) := x"07e0";
    tmp(34067) := x"07e0";
    tmp(34068) := x"07e0";
    tmp(34069) := x"07e0";
    tmp(34070) := x"07e0";
    tmp(34071) := x"07e0";
    tmp(34072) := x"07e0";
    tmp(34073) := x"07e0";
    tmp(34074) := x"07e0";
    tmp(34075) := x"07e0";
    tmp(34076) := x"07e0";
    tmp(34077) := x"0840";
    tmp(34078) := x"0840";
    tmp(34079) := x"0840";
    tmp(34080) := x"0020";
    tmp(34081) := x"00e5";
    tmp(34082) := x"00a3";
    tmp(34083) := x"0082";
    tmp(34084) := x"00c4";
    tmp(34085) := x"00e5";
    tmp(34086) := x"0105";
    tmp(34087) := x"0105";
    tmp(34088) := x"0105";
    tmp(34089) := x"0105";
    tmp(34090) := x"0105";
    tmp(34091) := x"00e5";
    tmp(34092) := x"00c4";
    tmp(34093) := x"00e5";
    tmp(34094) := x"0105";
    tmp(34095) := x"0105";
    tmp(34096) := x"0105";
    tmp(34097) := x"0105";
    tmp(34098) := x"0105";
    tmp(34099) := x"0925";
    tmp(34100) := x"0925";
    tmp(34101) := x"0926";
    tmp(34102) := x"0925";
    tmp(34103) := x"08e4";
    tmp(34104) := x"08c3";
    tmp(34105) := x"08e4";
    tmp(34106) := x"08e5";
    tmp(34107) := x"08e4";
    tmp(34108) := x"0905";
    tmp(34109) := x"0905";
    tmp(34110) := x"0905";
    tmp(34111) := x"0926";
    tmp(34112) := x"0926";
    tmp(34113) := x"08e5";
    tmp(34114) := x"0926";
    tmp(34115) := x"0947";
    tmp(34116) := x"0968";
    tmp(34117) := x"0988";
    tmp(34118) := x"0967";
    tmp(34119) := x"0905";
    tmp(34120) := x"08e5";
    tmp(34121) := x"0926";
    tmp(34122) := x"0988";
    tmp(34123) := x"0966";
    tmp(34124) := x"11e9";
    tmp(34125) := x"120a";
    tmp(34126) := x"11c8";
    tmp(34127) := x"11e6";
    tmp(34128) := x"19e4";
    tmp(34129) := x"1141";
    tmp(34130) := x"1141";
    tmp(34131) := x"1140";
    tmp(34132) := x"1140";
    tmp(34133) := x"1140";
    tmp(34134) := x"1140";
    tmp(34135) := x"1141";
    tmp(34136) := x"1161";
    tmp(34137) := x"1161";
    tmp(34138) := x"1161";
    tmp(34139) := x"1161";
    tmp(34140) := x"1161";
    tmp(34141) := x"1141";
    tmp(34142) := x"1161";
    tmp(34143) := x"1141";
    tmp(34144) := x"1161";
    tmp(34145) := x"1140";
    tmp(34146) := x"1140";
    tmp(34147) := x"1140";
    tmp(34148) := x"1140";
    tmp(34149) := x"0920";
    tmp(34150) := x"0920";
    tmp(34151) := x"0900";
    tmp(34152) := x"0900";
    tmp(34153) := x"08e0";
    tmp(34154) := x"08e0";
    tmp(34155) := x"0900";
    tmp(34156) := x"0900";
    tmp(34157) := x"08e1";
    tmp(34158) := x"10e1";
    tmp(34159) := x"1101";
    tmp(34160) := x"1101";
    tmp(34161) := x"1101";
    tmp(34162) := x"1102";
    tmp(34163) := x"1102";
    tmp(34164) := x"1902";
    tmp(34165) := x"1902";
    tmp(34166) := x"1902";
    tmp(34167) := x"1902";
    tmp(34168) := x"1902";
    tmp(34169) := x"1922";
    tmp(34170) := x"2123";
    tmp(34171) := x"1903";
    tmp(34172) := x"2102";
    tmp(34173) := x"2123";
    tmp(34174) := x"2143";
    tmp(34175) := x"2943";
    tmp(34176) := x"2964";
    tmp(34177) := x"2983";
    tmp(34178) := x"2983";
    tmp(34179) := x"2143";
    tmp(34180) := x"2142";
    tmp(34181) := x"1942";
    tmp(34182) := x"1942";
    tmp(34183) := x"1941";
    tmp(34184) := x"1921";
    tmp(34185) := x"1921";
    tmp(34186) := x"1921";
    tmp(34187) := x"1121";
    tmp(34188) := x"1121";
    tmp(34189) := x"1121";
    tmp(34190) := x"1101";
    tmp(34191) := x"0900";
    tmp(34192) := x"0900";
    tmp(34193) := x"0900";
    tmp(34194) := x"0900";
    tmp(34195) := x"1100";
    tmp(34196) := x"1100";
    tmp(34197) := x"1100";
    tmp(34198) := x"1100";
    tmp(34199) := x"1120";
    tmp(34200) := x"1100";
    tmp(34201) := x"10e0";
    tmp(34202) := x"1100";
    tmp(34203) := x"1100";
    tmp(34204) := x"1120";
    tmp(34205) := x"1121";
    tmp(34206) := x"1141";
    tmp(34207) := x"1120";
    tmp(34208) := x"1140";
    tmp(34209) := x"1120";
    tmp(34210) := x"0920";
    tmp(34211) := x"0920";
    tmp(34212) := x"0920";
    tmp(34213) := x"0900";
    tmp(34214) := x"0920";
    tmp(34215) := x"0900";
    tmp(34216) := x"1100";
    tmp(34217) := x"1100";
    tmp(34218) := x"10e0";
    tmp(34219) := x"1100";
    tmp(34220) := x"1100";
    tmp(34221) := x"1100";
    tmp(34222) := x"1100";
    tmp(34223) := x"10e0";
    tmp(34224) := x"10e0";
    tmp(34225) := x"10e0";
    tmp(34226) := x"18e0";
    tmp(34227) := x"18e1";
    tmp(34228) := x"18e1";
    tmp(34229) := x"18e1";
    tmp(34230) := x"18e1";
    tmp(34231) := x"18e1";
    tmp(34232) := x"10c1";
    tmp(34233) := x"10c1";
    tmp(34234) := x"10a1";
    tmp(34235) := x"10a0";
    tmp(34236) := x"1080";
    tmp(34237) := x"1080";
    tmp(34238) := x"0880";
    tmp(34239) := x"1060";
    tmp(34240) := x"1060";
    tmp(34241) := x"0860";
    tmp(34242) := x"0860";
    tmp(34243) := x"1060";
    tmp(34244) := x"1080";
    tmp(34245) := x"1080";
    tmp(34246) := x"1080";
    tmp(34247) := x"1080";
    tmp(34248) := x"1080";
    tmp(34249) := x"1080";
    tmp(34250) := x"1080";
    tmp(34251) := x"1081";
    tmp(34252) := x"1061";
    tmp(34253) := x"1061";
    tmp(34254) := x"1061";
    tmp(34255) := x"1061";
    tmp(34256) := x"1061";
    tmp(34257) := x"1061";
    tmp(34258) := x"1061";
    tmp(34259) := x"1061";
    tmp(34260) := x"1061";
    tmp(34261) := x"1061";
    tmp(34262) := x"1061";
    tmp(34263) := x"1061";
    tmp(34264) := x"1061";
    tmp(34265) := x"1060";
    tmp(34266) := x"1040";
    tmp(34267) := x"1060";
    tmp(34268) := x"1040";
    tmp(34269) := x"1040";
    tmp(34270) := x"1040";
    tmp(34271) := x"1040";
    tmp(34272) := x"1040";
    tmp(34273) := x"1040";
    tmp(34274) := x"1040";
    tmp(34275) := x"0840";
    tmp(34276) := x"0840";
    tmp(34277) := x"07e0";
    tmp(34278) := x"07e0";
    tmp(34279) := x"07e0";
    tmp(34280) := x"07e0";
    tmp(34281) := x"07e0";
    tmp(34282) := x"07e0";
    tmp(34283) := x"07e0";
    tmp(34284) := x"07e0";
    tmp(34285) := x"07e0";
    tmp(34286) := x"07e0";
    tmp(34287) := x"07e0";
    tmp(34288) := x"07e0";
    tmp(34289) := x"07e0";
    tmp(34290) := x"07e0";
    tmp(34291) := x"07e0";
    tmp(34292) := x"07e0";
    tmp(34293) := x"07e0";
    tmp(34294) := x"07e0";
    tmp(34295) := x"07e0";
    tmp(34296) := x"07e0";
    tmp(34297) := x"07e0";
    tmp(34298) := x"07e0";
    tmp(34299) := x"07e0";
    tmp(34300) := x"07e0";
    tmp(34301) := x"07e0";
    tmp(34302) := x"07e0";
    tmp(34303) := x"07e0";
    tmp(34304) := x"07e0";
    tmp(34305) := x"07e0";
    tmp(34306) := x"07e0";
    tmp(34307) := x"07e0";
    tmp(34308) := x"07e0";
    tmp(34309) := x"07e0";
    tmp(34310) := x"07e0";
    tmp(34311) := x"07e0";
    tmp(34312) := x"07e0";
    tmp(34313) := x"07e0";
    tmp(34314) := x"07e0";
    tmp(34315) := x"07e0";
    tmp(34316) := x"07e0";
    tmp(34317) := x"0840";
    tmp(34318) := x"0840";
    tmp(34319) := x"0840";
    tmp(34320) := x"0020";
    tmp(34321) := x"00e5";
    tmp(34322) := x"00a3";
    tmp(34323) := x"00a3";
    tmp(34324) := x"00e5";
    tmp(34325) := x"0105";
    tmp(34326) := x"0126";
    tmp(34327) := x"0126";
    tmp(34328) := x"0926";
    tmp(34329) := x"0125";
    tmp(34330) := x"0105";
    tmp(34331) := x"00e5";
    tmp(34332) := x"00e5";
    tmp(34333) := x"0105";
    tmp(34334) := x"0125";
    tmp(34335) := x"0126";
    tmp(34336) := x"0926";
    tmp(34337) := x"0126";
    tmp(34338) := x"0926";
    tmp(34339) := x"0946";
    tmp(34340) := x"0946";
    tmp(34341) := x"0925";
    tmp(34342) := x"00c3";
    tmp(34343) := x"08a3";
    tmp(34344) := x"08e4";
    tmp(34345) := x"0926";
    tmp(34346) := x"0926";
    tmp(34347) := x"0925";
    tmp(34348) := x"08e5";
    tmp(34349) := x"0905";
    tmp(34350) := x"0926";
    tmp(34351) := x"0925";
    tmp(34352) := x"0926";
    tmp(34353) := x"0967";
    tmp(34354) := x"0967";
    tmp(34355) := x"09a9";
    tmp(34356) := x"09c9";
    tmp(34357) := x"09c9";
    tmp(34358) := x"0946";
    tmp(34359) := x"0926";
    tmp(34360) := x"0926";
    tmp(34361) := x"09a8";
    tmp(34362) := x"122b";
    tmp(34363) := x"11a8";
    tmp(34364) := x"122a";
    tmp(34365) := x"1187";
    tmp(34366) := x"0944";
    tmp(34367) := x"1a03";
    tmp(34368) := x"1161";
    tmp(34369) := x"1141";
    tmp(34370) := x"1161";
    tmp(34371) := x"1161";
    tmp(34372) := x"1141";
    tmp(34373) := x"1141";
    tmp(34374) := x"1141";
    tmp(34375) := x"1141";
    tmp(34376) := x"1161";
    tmp(34377) := x"1161";
    tmp(34378) := x"1161";
    tmp(34379) := x"1161";
    tmp(34380) := x"1161";
    tmp(34381) := x"1141";
    tmp(34382) := x"1161";
    tmp(34383) := x"1141";
    tmp(34384) := x"1140";
    tmp(34385) := x"1140";
    tmp(34386) := x"1120";
    tmp(34387) := x"1120";
    tmp(34388) := x"1120";
    tmp(34389) := x"0920";
    tmp(34390) := x"0900";
    tmp(34391) := x"0900";
    tmp(34392) := x"0900";
    tmp(34393) := x"08e0";
    tmp(34394) := x"08e0";
    tmp(34395) := x"0900";
    tmp(34396) := x"08e0";
    tmp(34397) := x"0901";
    tmp(34398) := x"08e1";
    tmp(34399) := x"1101";
    tmp(34400) := x"1101";
    tmp(34401) := x"1101";
    tmp(34402) := x"1101";
    tmp(34403) := x"1102";
    tmp(34404) := x"1102";
    tmp(34405) := x"1902";
    tmp(34406) := x"1902";
    tmp(34407) := x"1902";
    tmp(34408) := x"1902";
    tmp(34409) := x"1902";
    tmp(34410) := x"1922";
    tmp(34411) := x"1902";
    tmp(34412) := x"1902";
    tmp(34413) := x"2123";
    tmp(34414) := x"2143";
    tmp(34415) := x"2943";
    tmp(34416) := x"2943";
    tmp(34417) := x"2943";
    tmp(34418) := x"2142";
    tmp(34419) := x"2142";
    tmp(34420) := x"1922";
    tmp(34421) := x"1921";
    tmp(34422) := x"1921";
    tmp(34423) := x"1921";
    tmp(34424) := x"1921";
    tmp(34425) := x"1121";
    tmp(34426) := x"1121";
    tmp(34427) := x"1121";
    tmp(34428) := x"1101";
    tmp(34429) := x"1101";
    tmp(34430) := x"0921";
    tmp(34431) := x"0900";
    tmp(34432) := x"0900";
    tmp(34433) := x"0900";
    tmp(34434) := x"1100";
    tmp(34435) := x"1100";
    tmp(34436) := x"1100";
    tmp(34437) := x"1100";
    tmp(34438) := x"1120";
    tmp(34439) := x"1100";
    tmp(34440) := x"1100";
    tmp(34441) := x"1100";
    tmp(34442) := x"1100";
    tmp(34443) := x"1100";
    tmp(34444) := x"1100";
    tmp(34445) := x"1121";
    tmp(34446) := x"1941";
    tmp(34447) := x"1120";
    tmp(34448) := x"1140";
    tmp(34449) := x"1120";
    tmp(34450) := x"0900";
    tmp(34451) := x"0920";
    tmp(34452) := x"0920";
    tmp(34453) := x"0920";
    tmp(34454) := x"0920";
    tmp(34455) := x"0900";
    tmp(34456) := x"0900";
    tmp(34457) := x"1100";
    tmp(34458) := x"1100";
    tmp(34459) := x"10e0";
    tmp(34460) := x"1100";
    tmp(34461) := x"10e0";
    tmp(34462) := x"10e0";
    tmp(34463) := x"10e0";
    tmp(34464) := x"10e0";
    tmp(34465) := x"10e0";
    tmp(34466) := x"10e0";
    tmp(34467) := x"18e0";
    tmp(34468) := x"18e0";
    tmp(34469) := x"18c1";
    tmp(34470) := x"18c0";
    tmp(34471) := x"10c0";
    tmp(34472) := x"10c1";
    tmp(34473) := x"10a0";
    tmp(34474) := x"10a0";
    tmp(34475) := x"10a0";
    tmp(34476) := x"0880";
    tmp(34477) := x"0880";
    tmp(34478) := x"0860";
    tmp(34479) := x"0860";
    tmp(34480) := x"0860";
    tmp(34481) := x"0860";
    tmp(34482) := x"1060";
    tmp(34483) := x"0860";
    tmp(34484) := x"1060";
    tmp(34485) := x"1080";
    tmp(34486) := x"1060";
    tmp(34487) := x"1080";
    tmp(34488) := x"1060";
    tmp(34489) := x"1080";
    tmp(34490) := x"1080";
    tmp(34491) := x"1060";
    tmp(34492) := x"1060";
    tmp(34493) := x"1060";
    tmp(34494) := x"1060";
    tmp(34495) := x"1061";
    tmp(34496) := x"1061";
    tmp(34497) := x"1061";
    tmp(34498) := x"1061";
    tmp(34499) := x"1061";
    tmp(34500) := x"1060";
    tmp(34501) := x"1060";
    tmp(34502) := x"1060";
    tmp(34503) := x"1060";
    tmp(34504) := x"1040";
    tmp(34505) := x"1040";
    tmp(34506) := x"1060";
    tmp(34507) := x"1040";
    tmp(34508) := x"1040";
    tmp(34509) := x"1040";
    tmp(34510) := x"1040";
    tmp(34511) := x"1040";
    tmp(34512) := x"1040";
    tmp(34513) := x"0840";
    tmp(34514) := x"0840";
    tmp(34515) := x"0840";
    tmp(34516) := x"0840";
    tmp(34517) := x"07e0";
    tmp(34518) := x"07e0";
    tmp(34519) := x"07e0";
    tmp(34520) := x"07e0";
    tmp(34521) := x"07e0";
    tmp(34522) := x"07e0";
    tmp(34523) := x"07e0";
    tmp(34524) := x"07e0";
    tmp(34525) := x"07e0";
    tmp(34526) := x"07e0";
    tmp(34527) := x"07e0";
    tmp(34528) := x"07e0";
    tmp(34529) := x"07e0";
    tmp(34530) := x"07e0";
    tmp(34531) := x"07e0";
    tmp(34532) := x"07e0";
    tmp(34533) := x"07e0";
    tmp(34534) := x"07e0";
    tmp(34535) := x"07e0";
    tmp(34536) := x"07e0";
    tmp(34537) := x"07e0";
    tmp(34538) := x"07e0";
    tmp(34539) := x"07e0";
    tmp(34540) := x"07e0";
    tmp(34541) := x"07e0";
    tmp(34542) := x"07e0";
    tmp(34543) := x"07e0";
    tmp(34544) := x"07e0";
    tmp(34545) := x"07e0";
    tmp(34546) := x"07e0";
    tmp(34547) := x"07e0";
    tmp(34548) := x"07e0";
    tmp(34549) := x"07e0";
    tmp(34550) := x"07e0";
    tmp(34551) := x"07e0";
    tmp(34552) := x"07e0";
    tmp(34553) := x"07e0";
    tmp(34554) := x"07e0";
    tmp(34555) := x"07e0";
    tmp(34556) := x"07e0";
    tmp(34557) := x"0840";
    tmp(34558) := x"0840";
    tmp(34559) := x"0840";
    tmp(34560) := x"0020";
    tmp(34561) := x"00e5";
    tmp(34562) := x"00a4";
    tmp(34563) := x"00a4";
    tmp(34564) := x"00e4";
    tmp(34565) := x"0105";
    tmp(34566) := x"0105";
    tmp(34567) := x"0105";
    tmp(34568) := x"0105";
    tmp(34569) := x"0105";
    tmp(34570) := x"00e5";
    tmp(34571) := x"00e5";
    tmp(34572) := x"0105";
    tmp(34573) := x"0126";
    tmp(34574) := x"0105";
    tmp(34575) := x"0105";
    tmp(34576) := x"00e5";
    tmp(34577) := x"00e4";
    tmp(34578) := x"0105";
    tmp(34579) := x"0905";
    tmp(34580) := x"0905";
    tmp(34581) := x"0905";
    tmp(34582) := x"08e4";
    tmp(34583) := x"00c3";
    tmp(34584) := x"08c4";
    tmp(34585) := x"00a3";
    tmp(34586) := x"00c4";
    tmp(34587) := x"0905";
    tmp(34588) := x"0926";
    tmp(34589) := x"0946";
    tmp(34590) := x"0946";
    tmp(34591) := x"0946";
    tmp(34592) := x"0966";
    tmp(34593) := x"0967";
    tmp(34594) := x"0967";
    tmp(34595) := x"0947";
    tmp(34596) := x"0947";
    tmp(34597) := x"0947";
    tmp(34598) := x"0967";
    tmp(34599) := x"0946";
    tmp(34600) := x"11a9";
    tmp(34601) := x"122b";
    tmp(34602) := x"11ea";
    tmp(34603) := x"1aac";
    tmp(34604) := x"11c7";
    tmp(34605) := x"1164";
    tmp(34606) := x"19c3";
    tmp(34607) := x"1161";
    tmp(34608) := x"1161";
    tmp(34609) := x"1161";
    tmp(34610) := x"1161";
    tmp(34611) := x"1161";
    tmp(34612) := x"1141";
    tmp(34613) := x"1141";
    tmp(34614) := x"1140";
    tmp(34615) := x"1141";
    tmp(34616) := x"1140";
    tmp(34617) := x"1160";
    tmp(34618) := x"1160";
    tmp(34619) := x"1160";
    tmp(34620) := x"1161";
    tmp(34621) := x"1141";
    tmp(34622) := x"1161";
    tmp(34623) := x"1141";
    tmp(34624) := x"1160";
    tmp(34625) := x"1140";
    tmp(34626) := x"1120";
    tmp(34627) := x"1120";
    tmp(34628) := x"0920";
    tmp(34629) := x"0920";
    tmp(34630) := x"0900";
    tmp(34631) := x"0900";
    tmp(34632) := x"08e0";
    tmp(34633) := x"08e0";
    tmp(34634) := x"08e0";
    tmp(34635) := x"08e0";
    tmp(34636) := x"08e0";
    tmp(34637) := x"08e0";
    tmp(34638) := x"0901";
    tmp(34639) := x"08e1";
    tmp(34640) := x"1101";
    tmp(34641) := x"1101";
    tmp(34642) := x"1101";
    tmp(34643) := x"1101";
    tmp(34644) := x"1102";
    tmp(34645) := x"1102";
    tmp(34646) := x"1902";
    tmp(34647) := x"1902";
    tmp(34648) := x"1902";
    tmp(34649) := x"1902";
    tmp(34650) := x"1902";
    tmp(34651) := x"1902";
    tmp(34652) := x"1922";
    tmp(34653) := x"2122";
    tmp(34654) := x"2123";
    tmp(34655) := x"2123";
    tmp(34656) := x"2143";
    tmp(34657) := x"2122";
    tmp(34658) := x"2122";
    tmp(34659) := x"1922";
    tmp(34660) := x"1921";
    tmp(34661) := x"1921";
    tmp(34662) := x"1921";
    tmp(34663) := x"1921";
    tmp(34664) := x"1921";
    tmp(34665) := x"1921";
    tmp(34666) := x"1121";
    tmp(34667) := x"1121";
    tmp(34668) := x"1101";
    tmp(34669) := x"1101";
    tmp(34670) := x"0900";
    tmp(34671) := x"08e0";
    tmp(34672) := x"0900";
    tmp(34673) := x"1100";
    tmp(34674) := x"1100";
    tmp(34675) := x"10e0";
    tmp(34676) := x"1100";
    tmp(34677) := x"1100";
    tmp(34678) := x"1100";
    tmp(34679) := x"1100";
    tmp(34680) := x"1100";
    tmp(34681) := x"1100";
    tmp(34682) := x"1100";
    tmp(34683) := x"1100";
    tmp(34684) := x"1100";
    tmp(34685) := x"1141";
    tmp(34686) := x"1941";
    tmp(34687) := x"1141";
    tmp(34688) := x"1140";
    tmp(34689) := x"1120";
    tmp(34690) := x"0920";
    tmp(34691) := x"0920";
    tmp(34692) := x"0920";
    tmp(34693) := x"0900";
    tmp(34694) := x"0900";
    tmp(34695) := x"0900";
    tmp(34696) := x"0900";
    tmp(34697) := x"08e0";
    tmp(34698) := x"08e0";
    tmp(34699) := x"08e0";
    tmp(34700) := x"10e0";
    tmp(34701) := x"10e0";
    tmp(34702) := x"10e0";
    tmp(34703) := x"10e0";
    tmp(34704) := x"10e0";
    tmp(34705) := x"10e0";
    tmp(34706) := x"10c0";
    tmp(34707) := x"10e0";
    tmp(34708) := x"18c0";
    tmp(34709) := x"10c0";
    tmp(34710) := x"10c0";
    tmp(34711) := x"10a0";
    tmp(34712) := x"10a0";
    tmp(34713) := x"10a0";
    tmp(34714) := x"1080";
    tmp(34715) := x"0880";
    tmp(34716) := x"0880";
    tmp(34717) := x"0880";
    tmp(34718) := x"0860";
    tmp(34719) := x"0860";
    tmp(34720) := x"0860";
    tmp(34721) := x"0860";
    tmp(34722) := x"0860";
    tmp(34723) := x"1060";
    tmp(34724) := x"1060";
    tmp(34725) := x"1060";
    tmp(34726) := x"1060";
    tmp(34727) := x"1080";
    tmp(34728) := x"1080";
    tmp(34729) := x"1060";
    tmp(34730) := x"1060";
    tmp(34731) := x"1060";
    tmp(34732) := x"1060";
    tmp(34733) := x"1060";
    tmp(34734) := x"1060";
    tmp(34735) := x"1060";
    tmp(34736) := x"1060";
    tmp(34737) := x"1060";
    tmp(34738) := x"1061";
    tmp(34739) := x"1060";
    tmp(34740) := x"1060";
    tmp(34741) := x"1060";
    tmp(34742) := x"1040";
    tmp(34743) := x"1040";
    tmp(34744) := x"1040";
    tmp(34745) := x"1040";
    tmp(34746) := x"1040";
    tmp(34747) := x"1040";
    tmp(34748) := x"1040";
    tmp(34749) := x"1040";
    tmp(34750) := x"0840";
    tmp(34751) := x"0840";
    tmp(34752) := x"0840";
    tmp(34753) := x"0840";
    tmp(34754) := x"0840";
    tmp(34755) := x"0840";
    tmp(34756) := x"0840";
    tmp(34757) := x"07e0";
    tmp(34758) := x"07e0";
    tmp(34759) := x"07e0";
    tmp(34760) := x"07e0";
    tmp(34761) := x"07e0";
    tmp(34762) := x"07e0";
    tmp(34763) := x"07e0";
    tmp(34764) := x"07e0";
    tmp(34765) := x"07e0";
    tmp(34766) := x"07e0";
    tmp(34767) := x"07e0";
    tmp(34768) := x"07e0";
    tmp(34769) := x"07e0";
    tmp(34770) := x"07e0";
    tmp(34771) := x"07e0";
    tmp(34772) := x"07e0";
    tmp(34773) := x"07e0";
    tmp(34774) := x"07e0";
    tmp(34775) := x"07e0";
    tmp(34776) := x"07e0";
    tmp(34777) := x"07e0";
    tmp(34778) := x"07e0";
    tmp(34779) := x"07e0";
    tmp(34780) := x"07e0";
    tmp(34781) := x"07e0";
    tmp(34782) := x"07e0";
    tmp(34783) := x"07e0";
    tmp(34784) := x"07e0";
    tmp(34785) := x"07e0";
    tmp(34786) := x"07e0";
    tmp(34787) := x"07e0";
    tmp(34788) := x"07e0";
    tmp(34789) := x"07e0";
    tmp(34790) := x"07e0";
    tmp(34791) := x"07e0";
    tmp(34792) := x"07e0";
    tmp(34793) := x"07e0";
    tmp(34794) := x"07e0";
    tmp(34795) := x"07e0";
    tmp(34796) := x"07e0";
    tmp(34797) := x"0840";
    tmp(34798) := x"0840";
    tmp(34799) := x"0840";
    tmp(34800) := x"0020";
    tmp(34801) := x"00e5";
    tmp(34802) := x"0083";
    tmp(34803) := x"00c4";
    tmp(34804) := x"00e4";
    tmp(34805) := x"00e4";
    tmp(34806) := x"00e4";
    tmp(34807) := x"00e4";
    tmp(34808) := x"00e4";
    tmp(34809) := x"00e4";
    tmp(34810) := x"00c4";
    tmp(34811) := x"00c4";
    tmp(34812) := x"00e4";
    tmp(34813) := x"00c4";
    tmp(34814) := x"00c4";
    tmp(34815) := x"00e4";
    tmp(34816) := x"00e4";
    tmp(34817) := x"00e4";
    tmp(34818) := x"00e4";
    tmp(34819) := x"00e4";
    tmp(34820) := x"00e4";
    tmp(34821) := x"00e4";
    tmp(34822) := x"00e4";
    tmp(34823) := x"00c4";
    tmp(34824) := x"00c4";
    tmp(34825) := x"00c4";
    tmp(34826) := x"0926";
    tmp(34827) := x"0988";
    tmp(34828) := x"09a8";
    tmp(34829) := x"0967";
    tmp(34830) := x"0946";
    tmp(34831) := x"0946";
    tmp(34832) := x"0966";
    tmp(34833) := x"0926";
    tmp(34834) := x"0967";
    tmp(34835) := x"0988";
    tmp(34836) := x"09a8";
    tmp(34837) := x"11e9";
    tmp(34838) := x"09a7";
    tmp(34839) := x"0926";
    tmp(34840) := x"0987";
    tmp(34841) := x"0967";
    tmp(34842) := x"120a";
    tmp(34843) := x"0966";
    tmp(34844) := x"1164";
    tmp(34845) := x"1162";
    tmp(34846) := x"1161";
    tmp(34847) := x"1161";
    tmp(34848) := x"1161";
    tmp(34849) := x"1161";
    tmp(34850) := x"1161";
    tmp(34851) := x"1141";
    tmp(34852) := x"1140";
    tmp(34853) := x"1140";
    tmp(34854) := x"1140";
    tmp(34855) := x"1141";
    tmp(34856) := x"1140";
    tmp(34857) := x"1160";
    tmp(34858) := x"1140";
    tmp(34859) := x"1161";
    tmp(34860) := x"1161";
    tmp(34861) := x"1161";
    tmp(34862) := x"1161";
    tmp(34863) := x"1140";
    tmp(34864) := x"1140";
    tmp(34865) := x"1140";
    tmp(34866) := x"1140";
    tmp(34867) := x"0920";
    tmp(34868) := x"0920";
    tmp(34869) := x"0900";
    tmp(34870) := x"0900";
    tmp(34871) := x"0900";
    tmp(34872) := x"08e0";
    tmp(34873) := x"08e0";
    tmp(34874) := x"08e0";
    tmp(34875) := x"08e0";
    tmp(34876) := x"08e0";
    tmp(34877) := x"0900";
    tmp(34878) := x"0900";
    tmp(34879) := x"08e1";
    tmp(34880) := x"1101";
    tmp(34881) := x"10e1";
    tmp(34882) := x"1101";
    tmp(34883) := x"1101";
    tmp(34884) := x"1101";
    tmp(34885) := x"1102";
    tmp(34886) := x"1102";
    tmp(34887) := x"1902";
    tmp(34888) := x"1902";
    tmp(34889) := x"1902";
    tmp(34890) := x"1902";
    tmp(34891) := x"1902";
    tmp(34892) := x"1922";
    tmp(34893) := x"2122";
    tmp(34894) := x"2122";
    tmp(34895) := x"2122";
    tmp(34896) := x"2122";
    tmp(34897) := x"2122";
    tmp(34898) := x"1922";
    tmp(34899) := x"1921";
    tmp(34900) := x"1921";
    tmp(34901) := x"1921";
    tmp(34902) := x"1921";
    tmp(34903) := x"1921";
    tmp(34904) := x"1921";
    tmp(34905) := x"1121";
    tmp(34906) := x"1121";
    tmp(34907) := x"1101";
    tmp(34908) := x"1121";
    tmp(34909) := x"0900";
    tmp(34910) := x"0900";
    tmp(34911) := x"0900";
    tmp(34912) := x"1100";
    tmp(34913) := x"1100";
    tmp(34914) := x"1100";
    tmp(34915) := x"1100";
    tmp(34916) := x"1100";
    tmp(34917) := x"1100";
    tmp(34918) := x"1100";
    tmp(34919) := x"1100";
    tmp(34920) := x"1100";
    tmp(34921) := x"1100";
    tmp(34922) := x"1100";
    tmp(34923) := x"1100";
    tmp(34924) := x"1100";
    tmp(34925) := x"1121";
    tmp(34926) := x"1120";
    tmp(34927) := x"1141";
    tmp(34928) := x"1141";
    tmp(34929) := x"1120";
    tmp(34930) := x"0920";
    tmp(34931) := x"0900";
    tmp(34932) := x"0900";
    tmp(34933) := x"0920";
    tmp(34934) := x"0920";
    tmp(34935) := x"0900";
    tmp(34936) := x"0900";
    tmp(34937) := x"0900";
    tmp(34938) := x"08e0";
    tmp(34939) := x"08e0";
    tmp(34940) := x"08e0";
    tmp(34941) := x"10e0";
    tmp(34942) := x"10e0";
    tmp(34943) := x"10e0";
    tmp(34944) := x"10c0";
    tmp(34945) := x"10c0";
    tmp(34946) := x"10c0";
    tmp(34947) := x"10c0";
    tmp(34948) := x"10c0";
    tmp(34949) := x"10c0";
    tmp(34950) := x"10a0";
    tmp(34951) := x"10a0";
    tmp(34952) := x"10a0";
    tmp(34953) := x"1080";
    tmp(34954) := x"0880";
    tmp(34955) := x"0880";
    tmp(34956) := x"0880";
    tmp(34957) := x"0860";
    tmp(34958) := x"0860";
    tmp(34959) := x"0860";
    tmp(34960) := x"0860";
    tmp(34961) := x"1060";
    tmp(34962) := x"1060";
    tmp(34963) := x"1060";
    tmp(34964) := x"1060";
    tmp(34965) := x"1060";
    tmp(34966) := x"1060";
    tmp(34967) := x"1060";
    tmp(34968) := x"1060";
    tmp(34969) := x"1060";
    tmp(34970) := x"1060";
    tmp(34971) := x"1060";
    tmp(34972) := x"1060";
    tmp(34973) := x"1060";
    tmp(34974) := x"1040";
    tmp(34975) := x"1040";
    tmp(34976) := x"1040";
    tmp(34977) := x"1040";
    tmp(34978) := x"1040";
    tmp(34979) := x"1040";
    tmp(34980) := x"1060";
    tmp(34981) := x"1040";
    tmp(34982) := x"1040";
    tmp(34983) := x"1040";
    tmp(34984) := x"1040";
    tmp(34985) := x"1040";
    tmp(34986) := x"1040";
    tmp(34987) := x"1040";
    tmp(34988) := x"1040";
    tmp(34989) := x"1040";
    tmp(34990) := x"0840";
    tmp(34991) := x"0840";
    tmp(34992) := x"0840";
    tmp(34993) := x"0840";
    tmp(34994) := x"0840";
    tmp(34995) := x"0840";
    tmp(34996) := x"0840";
    tmp(34997) := x"07e0";
    tmp(34998) := x"07e0";
    tmp(34999) := x"07e0";
    tmp(35000) := x"07e0";
    tmp(35001) := x"07e0";
    tmp(35002) := x"07e0";
    tmp(35003) := x"07e0";
    tmp(35004) := x"07e0";
    tmp(35005) := x"07e0";
    tmp(35006) := x"07e0";
    tmp(35007) := x"07e0";
    tmp(35008) := x"07e0";
    tmp(35009) := x"07e0";
    tmp(35010) := x"07e0";
    tmp(35011) := x"07e0";
    tmp(35012) := x"07e0";
    tmp(35013) := x"07e0";
    tmp(35014) := x"07e0";
    tmp(35015) := x"07e0";
    tmp(35016) := x"07e0";
    tmp(35017) := x"07e0";
    tmp(35018) := x"07e0";
    tmp(35019) := x"07e0";
    tmp(35020) := x"07e0";
    tmp(35021) := x"07e0";
    tmp(35022) := x"07e0";
    tmp(35023) := x"07e0";
    tmp(35024) := x"07e0";
    tmp(35025) := x"07e0";
    tmp(35026) := x"07e0";
    tmp(35027) := x"07e0";
    tmp(35028) := x"07e0";
    tmp(35029) := x"07e0";
    tmp(35030) := x"07e0";
    tmp(35031) := x"07e0";
    tmp(35032) := x"07e0";
    tmp(35033) := x"07e0";
    tmp(35034) := x"07e0";
    tmp(35035) := x"07e0";
    tmp(35036) := x"07e0";
    tmp(35037) := x"0840";
    tmp(35038) := x"0840";
    tmp(35039) := x"0840";
    tmp(35040) := x"0020";
    tmp(35041) := x"00e4";
    tmp(35042) := x"00a3";
    tmp(35043) := x"00c4";
    tmp(35044) := x"00e4";
    tmp(35045) := x"00e5";
    tmp(35046) := x"00e5";
    tmp(35047) := x"00e4";
    tmp(35048) := x"00c4";
    tmp(35049) := x"00c4";
    tmp(35050) := x"00c3";
    tmp(35051) := x"00a3";
    tmp(35052) := x"00e5";
    tmp(35053) := x"00e5";
    tmp(35054) := x"0105";
    tmp(35055) := x"0105";
    tmp(35056) := x"0105";
    tmp(35057) := x"0105";
    tmp(35058) := x"00e5";
    tmp(35059) := x"0104";
    tmp(35060) := x"0905";
    tmp(35061) := x"00e4";
    tmp(35062) := x"00c4";
    tmp(35063) := x"0905";
    tmp(35064) := x"0926";
    tmp(35065) := x"0926";
    tmp(35066) := x"0947";
    tmp(35067) := x"0947";
    tmp(35068) := x"0947";
    tmp(35069) := x"0947";
    tmp(35070) := x"0967";
    tmp(35071) := x"0925";
    tmp(35072) := x"0924";
    tmp(35073) := x"0925";
    tmp(35074) := x"09a8";
    tmp(35075) := x"11ea";
    tmp(35076) := x"0988";
    tmp(35077) := x"0925";
    tmp(35078) := x"0966";
    tmp(35079) := x"1209";
    tmp(35080) := x"0925";
    tmp(35081) := x"0925";
    tmp(35082) := x"0966";
    tmp(35083) := x"11a5";
    tmp(35084) := x"0901";
    tmp(35085) := x"1161";
    tmp(35086) := x"1181";
    tmp(35087) := x"1141";
    tmp(35088) := x"1161";
    tmp(35089) := x"1161";
    tmp(35090) := x"1161";
    tmp(35091) := x"1140";
    tmp(35092) := x"1140";
    tmp(35093) := x"1140";
    tmp(35094) := x"1140";
    tmp(35095) := x"1160";
    tmp(35096) := x"1140";
    tmp(35097) := x"1140";
    tmp(35098) := x"1140";
    tmp(35099) := x"1160";
    tmp(35100) := x"1140";
    tmp(35101) := x"1141";
    tmp(35102) := x"1160";
    tmp(35103) := x"1140";
    tmp(35104) := x"1140";
    tmp(35105) := x"1140";
    tmp(35106) := x"1120";
    tmp(35107) := x"0920";
    tmp(35108) := x"0900";
    tmp(35109) := x"0900";
    tmp(35110) := x"0900";
    tmp(35111) := x"0900";
    tmp(35112) := x"08e0";
    tmp(35113) := x"08e0";
    tmp(35114) := x"08e0";
    tmp(35115) := x"08e0";
    tmp(35116) := x"08e0";
    tmp(35117) := x"0900";
    tmp(35118) := x"08e0";
    tmp(35119) := x"0901";
    tmp(35120) := x"08e1";
    tmp(35121) := x"1101";
    tmp(35122) := x"1101";
    tmp(35123) := x"1101";
    tmp(35124) := x"1102";
    tmp(35125) := x"1102";
    tmp(35126) := x"1102";
    tmp(35127) := x"1102";
    tmp(35128) := x"1902";
    tmp(35129) := x"1902";
    tmp(35130) := x"18e2";
    tmp(35131) := x"1902";
    tmp(35132) := x"1922";
    tmp(35133) := x"1902";
    tmp(35134) := x"1902";
    tmp(35135) := x"2122";
    tmp(35136) := x"2122";
    tmp(35137) := x"2122";
    tmp(35138) := x"1922";
    tmp(35139) := x"1921";
    tmp(35140) := x"1921";
    tmp(35141) := x"1901";
    tmp(35142) := x"1921";
    tmp(35143) := x"1941";
    tmp(35144) := x"1121";
    tmp(35145) := x"1121";
    tmp(35146) := x"1121";
    tmp(35147) := x"1101";
    tmp(35148) := x"1100";
    tmp(35149) := x"0900";
    tmp(35150) := x"08e0";
    tmp(35151) := x"08e0";
    tmp(35152) := x"1100";
    tmp(35153) := x"1100";
    tmp(35154) := x"1100";
    tmp(35155) := x"1100";
    tmp(35156) := x"10e0";
    tmp(35157) := x"1100";
    tmp(35158) := x"1100";
    tmp(35159) := x"1100";
    tmp(35160) := x"1100";
    tmp(35161) := x"1100";
    tmp(35162) := x"1100";
    tmp(35163) := x"1100";
    tmp(35164) := x"1121";
    tmp(35165) := x"1121";
    tmp(35166) := x"1120";
    tmp(35167) := x"1141";
    tmp(35168) := x"1141";
    tmp(35169) := x"1120";
    tmp(35170) := x"0920";
    tmp(35171) := x"0900";
    tmp(35172) := x"0920";
    tmp(35173) := x"0920";
    tmp(35174) := x"0900";
    tmp(35175) := x"0900";
    tmp(35176) := x"0900";
    tmp(35177) := x"0900";
    tmp(35178) := x"08e0";
    tmp(35179) := x"08e0";
    tmp(35180) := x"08e0";
    tmp(35181) := x"08e0";
    tmp(35182) := x"10c0";
    tmp(35183) := x"10c0";
    tmp(35184) := x"10c0";
    tmp(35185) := x"10c0";
    tmp(35186) := x"10c0";
    tmp(35187) := x"10c0";
    tmp(35188) := x"10c0";
    tmp(35189) := x"10a0";
    tmp(35190) := x"10a0";
    tmp(35191) := x"10a0";
    tmp(35192) := x"10a0";
    tmp(35193) := x"1080";
    tmp(35194) := x"1080";
    tmp(35195) := x"0860";
    tmp(35196) := x"0860";
    tmp(35197) := x"0860";
    tmp(35198) := x"0860";
    tmp(35199) := x"1060";
    tmp(35200) := x"1060";
    tmp(35201) := x"0860";
    tmp(35202) := x"1060";
    tmp(35203) := x"1060";
    tmp(35204) := x"1060";
    tmp(35205) := x"1060";
    tmp(35206) := x"1060";
    tmp(35207) := x"1060";
    tmp(35208) := x"1060";
    tmp(35209) := x"1060";
    tmp(35210) := x"1060";
    tmp(35211) := x"1060";
    tmp(35212) := x"1040";
    tmp(35213) := x"1040";
    tmp(35214) := x"1040";
    tmp(35215) := x"1040";
    tmp(35216) := x"1040";
    tmp(35217) := x"1040";
    tmp(35218) := x"1040";
    tmp(35219) := x"1040";
    tmp(35220) := x"1040";
    tmp(35221) := x"1060";
    tmp(35222) := x"1040";
    tmp(35223) := x"1040";
    tmp(35224) := x"1040";
    tmp(35225) := x"1040";
    tmp(35226) := x"1040";
    tmp(35227) := x"1040";
    tmp(35228) := x"1040";
    tmp(35229) := x"1040";
    tmp(35230) := x"1040";
    tmp(35231) := x"0840";
    tmp(35232) := x"0840";
    tmp(35233) := x"0840";
    tmp(35234) := x"0840";
    tmp(35235) := x"0840";
    tmp(35236) := x"0840";
    tmp(35237) := x"07e0";
    tmp(35238) := x"07e0";
    tmp(35239) := x"07e0";
    tmp(35240) := x"07e0";
    tmp(35241) := x"07e0";
    tmp(35242) := x"07e0";
    tmp(35243) := x"07e0";
    tmp(35244) := x"07e0";
    tmp(35245) := x"07e0";
    tmp(35246) := x"07e0";
    tmp(35247) := x"07e0";
    tmp(35248) := x"07e0";
    tmp(35249) := x"07e0";
    tmp(35250) := x"07e0";
    tmp(35251) := x"07e0";
    tmp(35252) := x"07e0";
    tmp(35253) := x"07e0";
    tmp(35254) := x"07e0";
    tmp(35255) := x"07e0";
    tmp(35256) := x"07e0";
    tmp(35257) := x"07e0";
    tmp(35258) := x"07e0";
    tmp(35259) := x"07e0";
    tmp(35260) := x"07e0";
    tmp(35261) := x"07e0";
    tmp(35262) := x"07e0";
    tmp(35263) := x"07e0";
    tmp(35264) := x"07e0";
    tmp(35265) := x"07e0";
    tmp(35266) := x"07e0";
    tmp(35267) := x"07e0";
    tmp(35268) := x"07e0";
    tmp(35269) := x"07e0";
    tmp(35270) := x"07e0";
    tmp(35271) := x"07e0";
    tmp(35272) := x"07e0";
    tmp(35273) := x"07e0";
    tmp(35274) := x"07e0";
    tmp(35275) := x"07e0";
    tmp(35276) := x"07e0";
    tmp(35277) := x"0840";
    tmp(35278) := x"0840";
    tmp(35279) := x"0840";
    tmp(35280) := x"0020";
    tmp(35281) := x"00c4";
    tmp(35282) := x"00c4";
    tmp(35283) := x"0062";
    tmp(35284) := x"00a3";
    tmp(35285) := x"0105";
    tmp(35286) := x"0105";
    tmp(35287) := x"00e5";
    tmp(35288) := x"00c4";
    tmp(35289) := x"00c4";
    tmp(35290) := x"00c4";
    tmp(35291) := x"00c4";
    tmp(35292) := x"00c4";
    tmp(35293) := x"0105";
    tmp(35294) := x"0126";
    tmp(35295) := x"0126";
    tmp(35296) := x"0926";
    tmp(35297) := x"0926";
    tmp(35298) := x"0926";
    tmp(35299) := x"0926";
    tmp(35300) := x"0926";
    tmp(35301) := x"0925";
    tmp(35302) := x"0905";
    tmp(35303) := x"0906";
    tmp(35304) := x"0926";
    tmp(35305) := x"0946";
    tmp(35306) := x"0987";
    tmp(35307) := x"0987";
    tmp(35308) := x"0987";
    tmp(35309) := x"09a7";
    tmp(35310) := x"09a7";
    tmp(35311) := x"11a7";
    tmp(35312) := x"0986";
    tmp(35313) := x"0946";
    tmp(35314) := x"0905";
    tmp(35315) := x"00c4";
    tmp(35316) := x"0905";
    tmp(35317) := x"09c9";
    tmp(35318) := x"120a";
    tmp(35319) := x"0904";
    tmp(35320) := x"08c3";
    tmp(35321) := x"11a6";
    tmp(35322) := x"1164";
    tmp(35323) := x"0901";
    tmp(35324) := x"1161";
    tmp(35325) := x"1181";
    tmp(35326) := x"1161";
    tmp(35327) := x"1161";
    tmp(35328) := x"1161";
    tmp(35329) := x"1161";
    tmp(35330) := x"1140";
    tmp(35331) := x"1140";
    tmp(35332) := x"1140";
    tmp(35333) := x"1140";
    tmp(35334) := x"1140";
    tmp(35335) := x"1140";
    tmp(35336) := x"1140";
    tmp(35337) := x"1140";
    tmp(35338) := x"1140";
    tmp(35339) := x"1140";
    tmp(35340) := x"1140";
    tmp(35341) := x"1140";
    tmp(35342) := x"1140";
    tmp(35343) := x"1140";
    tmp(35344) := x"1140";
    tmp(35345) := x"1120";
    tmp(35346) := x"1120";
    tmp(35347) := x"0920";
    tmp(35348) := x"0920";
    tmp(35349) := x"0900";
    tmp(35350) := x"0900";
    tmp(35351) := x"0900";
    tmp(35352) := x"0900";
    tmp(35353) := x"0900";
    tmp(35354) := x"0900";
    tmp(35355) := x"08e0";
    tmp(35356) := x"08e0";
    tmp(35357) := x"0900";
    tmp(35358) := x"0900";
    tmp(35359) := x"0901";
    tmp(35360) := x"1101";
    tmp(35361) := x"1101";
    tmp(35362) := x"1101";
    tmp(35363) := x"1101";
    tmp(35364) := x"1101";
    tmp(35365) := x"1101";
    tmp(35366) := x"1102";
    tmp(35367) := x"1102";
    tmp(35368) := x"1102";
    tmp(35369) := x"1902";
    tmp(35370) := x"1922";
    tmp(35371) := x"1902";
    tmp(35372) := x"1902";
    tmp(35373) := x"1922";
    tmp(35374) := x"2122";
    tmp(35375) := x"2122";
    tmp(35376) := x"1922";
    tmp(35377) := x"1922";
    tmp(35378) := x"1921";
    tmp(35379) := x"1921";
    tmp(35380) := x"1921";
    tmp(35381) := x"1921";
    tmp(35382) := x"1921";
    tmp(35383) := x"1941";
    tmp(35384) := x"1121";
    tmp(35385) := x"1121";
    tmp(35386) := x"1101";
    tmp(35387) := x"1101";
    tmp(35388) := x"0900";
    tmp(35389) := x"0900";
    tmp(35390) := x"0900";
    tmp(35391) := x"0900";
    tmp(35392) := x"1100";
    tmp(35393) := x"1100";
    tmp(35394) := x"1100";
    tmp(35395) := x"1100";
    tmp(35396) := x"10e0";
    tmp(35397) := x"10e0";
    tmp(35398) := x"1100";
    tmp(35399) := x"1100";
    tmp(35400) := x"1100";
    tmp(35401) := x"1100";
    tmp(35402) := x"10e0";
    tmp(35403) := x"1100";
    tmp(35404) := x"1120";
    tmp(35405) := x"1120";
    tmp(35406) := x"1100";
    tmp(35407) := x"1120";
    tmp(35408) := x"1140";
    tmp(35409) := x"1140";
    tmp(35410) := x"0920";
    tmp(35411) := x"0900";
    tmp(35412) := x"0920";
    tmp(35413) := x"0920";
    tmp(35414) := x"0920";
    tmp(35415) := x"0900";
    tmp(35416) := x"0900";
    tmp(35417) := x"0900";
    tmp(35418) := x"08e0";
    tmp(35419) := x"08e0";
    tmp(35420) := x"08e0";
    tmp(35421) := x"08c0";
    tmp(35422) := x"08c0";
    tmp(35423) := x"08c0";
    tmp(35424) := x"08c0";
    tmp(35425) := x"10c0";
    tmp(35426) := x"10a0";
    tmp(35427) := x"10a0";
    tmp(35428) := x"10a0";
    tmp(35429) := x"10a0";
    tmp(35430) := x"10a0";
    tmp(35431) := x"1080";
    tmp(35432) := x"1080";
    tmp(35433) := x"0880";
    tmp(35434) := x"0880";
    tmp(35435) := x"0880";
    tmp(35436) := x"0860";
    tmp(35437) := x"0860";
    tmp(35438) := x"0860";
    tmp(35439) := x"0860";
    tmp(35440) := x"1060";
    tmp(35441) := x"1060";
    tmp(35442) := x"1060";
    tmp(35443) := x"1060";
    tmp(35444) := x"1060";
    tmp(35445) := x"1060";
    tmp(35446) := x"1060";
    tmp(35447) := x"1060";
    tmp(35448) := x"1060";
    tmp(35449) := x"1060";
    tmp(35450) := x"1060";
    tmp(35451) := x"1040";
    tmp(35452) := x"1040";
    tmp(35453) := x"1040";
    tmp(35454) := x"0840";
    tmp(35455) := x"1040";
    tmp(35456) := x"1040";
    tmp(35457) := x"1040";
    tmp(35458) := x"1040";
    tmp(35459) := x"1040";
    tmp(35460) := x"1040";
    tmp(35461) := x"1040";
    tmp(35462) := x"1040";
    tmp(35463) := x"1040";
    tmp(35464) := x"1040";
    tmp(35465) := x"1040";
    tmp(35466) := x"1040";
    tmp(35467) := x"1040";
    tmp(35468) := x"1040";
    tmp(35469) := x"1040";
    tmp(35470) := x"0840";
    tmp(35471) := x"0840";
    tmp(35472) := x"0840";
    tmp(35473) := x"1040";
    tmp(35474) := x"0840";
    tmp(35475) := x"0840";
    tmp(35476) := x"0840";
    tmp(35477) := x"07e0";
    tmp(35478) := x"07e0";
    tmp(35479) := x"07e0";
    tmp(35480) := x"07e0";
    tmp(35481) := x"07e0";
    tmp(35482) := x"07e0";
    tmp(35483) := x"07e0";
    tmp(35484) := x"07e0";
    tmp(35485) := x"07e0";
    tmp(35486) := x"07e0";
    tmp(35487) := x"07e0";
    tmp(35488) := x"07e0";
    tmp(35489) := x"07e0";
    tmp(35490) := x"07e0";
    tmp(35491) := x"07e0";
    tmp(35492) := x"07e0";
    tmp(35493) := x"07e0";
    tmp(35494) := x"07e0";
    tmp(35495) := x"07e0";
    tmp(35496) := x"07e0";
    tmp(35497) := x"07e0";
    tmp(35498) := x"07e0";
    tmp(35499) := x"07e0";
    tmp(35500) := x"07e0";
    tmp(35501) := x"07e0";
    tmp(35502) := x"07e0";
    tmp(35503) := x"07e0";
    tmp(35504) := x"07e0";
    tmp(35505) := x"07e0";
    tmp(35506) := x"07e0";
    tmp(35507) := x"07e0";
    tmp(35508) := x"07e0";
    tmp(35509) := x"07e0";
    tmp(35510) := x"07e0";
    tmp(35511) := x"07e0";
    tmp(35512) := x"07e0";
    tmp(35513) := x"07e0";
    tmp(35514) := x"07e0";
    tmp(35515) := x"07e0";
    tmp(35516) := x"07e0";
    tmp(35517) := x"0840";
    tmp(35518) := x"0840";
    tmp(35519) := x"0840";
    tmp(35520) := x"0020";
    tmp(35521) := x"00e5";
    tmp(35522) := x"00c4";
    tmp(35523) := x"0062";
    tmp(35524) := x"0082";
    tmp(35525) := x"00c4";
    tmp(35526) := x"0105";
    tmp(35527) := x"0106";
    tmp(35528) := x"00e5";
    tmp(35529) := x"00e5";
    tmp(35530) := x"00e5";
    tmp(35531) := x"00e4";
    tmp(35532) := x"00e4";
    tmp(35533) := x"00c4";
    tmp(35534) := x"00c4";
    tmp(35535) := x"00e5";
    tmp(35536) := x"0105";
    tmp(35537) := x"0926";
    tmp(35538) := x"0947";
    tmp(35539) := x"0968";
    tmp(35540) := x"0968";
    tmp(35541) := x"0947";
    tmp(35542) := x"0947";
    tmp(35543) := x"0967";
    tmp(35544) := x"09a9";
    tmp(35545) := x"09c9";
    tmp(35546) := x"09c9";
    tmp(35547) := x"09e9";
    tmp(35548) := x"11e9";
    tmp(35549) := x"120a";
    tmp(35550) := x"11e9";
    tmp(35551) := x"09a8";
    tmp(35552) := x"0925";
    tmp(35553) := x"0925";
    tmp(35554) := x"00e4";
    tmp(35555) := x"00a3";
    tmp(35556) := x"0967";
    tmp(35557) := x"0989";
    tmp(35558) := x"0926";
    tmp(35559) := x"0986";
    tmp(35560) := x"1185";
    tmp(35561) := x"08e2";
    tmp(35562) := x"1101";
    tmp(35563) := x"1981";
    tmp(35564) := x"1181";
    tmp(35565) := x"1161";
    tmp(35566) := x"1141";
    tmp(35567) := x"1140";
    tmp(35568) := x"1140";
    tmp(35569) := x"1140";
    tmp(35570) := x"1140";
    tmp(35571) := x"1140";
    tmp(35572) := x"1140";
    tmp(35573) := x"1120";
    tmp(35574) := x"1120";
    tmp(35575) := x"1140";
    tmp(35576) := x"1140";
    tmp(35577) := x"1140";
    tmp(35578) := x"1140";
    tmp(35579) := x"1120";
    tmp(35580) := x"1140";
    tmp(35581) := x"1140";
    tmp(35582) := x"1140";
    tmp(35583) := x"1140";
    tmp(35584) := x"1120";
    tmp(35585) := x"1120";
    tmp(35586) := x"0920";
    tmp(35587) := x"0920";
    tmp(35588) := x"0920";
    tmp(35589) := x"0920";
    tmp(35590) := x"0920";
    tmp(35591) := x"0920";
    tmp(35592) := x"0900";
    tmp(35593) := x"0900";
    tmp(35594) := x"0900";
    tmp(35595) := x"0900";
    tmp(35596) := x"08e0";
    tmp(35597) := x"0900";
    tmp(35598) := x"0900";
    tmp(35599) := x"0921";
    tmp(35600) := x"1101";
    tmp(35601) := x"1101";
    tmp(35602) := x"1101";
    tmp(35603) := x"1101";
    tmp(35604) := x"1121";
    tmp(35605) := x"1121";
    tmp(35606) := x"1122";
    tmp(35607) := x"1102";
    tmp(35608) := x"1102";
    tmp(35609) := x"1102";
    tmp(35610) := x"1902";
    tmp(35611) := x"1102";
    tmp(35612) := x"1902";
    tmp(35613) := x"1902";
    tmp(35614) := x"1922";
    tmp(35615) := x"1922";
    tmp(35616) := x"1921";
    tmp(35617) := x"1921";
    tmp(35618) := x"1921";
    tmp(35619) := x"1921";
    tmp(35620) := x"1921";
    tmp(35621) := x"1941";
    tmp(35622) := x"1921";
    tmp(35623) := x"1941";
    tmp(35624) := x"1121";
    tmp(35625) := x"1121";
    tmp(35626) := x"1101";
    tmp(35627) := x"1100";
    tmp(35628) := x"0900";
    tmp(35629) := x"08e0";
    tmp(35630) := x"08e0";
    tmp(35631) := x"1100";
    tmp(35632) := x"1100";
    tmp(35633) := x"1100";
    tmp(35634) := x"1100";
    tmp(35635) := x"1100";
    tmp(35636) := x"10e0";
    tmp(35637) := x"10e0";
    tmp(35638) := x"1100";
    tmp(35639) := x"1101";
    tmp(35640) := x"1101";
    tmp(35641) := x"1101";
    tmp(35642) := x"10e0";
    tmp(35643) := x"1100";
    tmp(35644) := x"1120";
    tmp(35645) := x"1100";
    tmp(35646) := x"1100";
    tmp(35647) := x"1120";
    tmp(35648) := x"1140";
    tmp(35649) := x"1140";
    tmp(35650) := x"1120";
    tmp(35651) := x"0900";
    tmp(35652) := x"0920";
    tmp(35653) := x"0900";
    tmp(35654) := x"0920";
    tmp(35655) := x"0900";
    tmp(35656) := x"0900";
    tmp(35657) := x"0900";
    tmp(35658) := x"08e0";
    tmp(35659) := x"08e0";
    tmp(35660) := x"08c0";
    tmp(35661) := x"08c0";
    tmp(35662) := x"08c0";
    tmp(35663) := x"08c0";
    tmp(35664) := x"08c0";
    tmp(35665) := x"10c0";
    tmp(35666) := x"08a0";
    tmp(35667) := x"10a0";
    tmp(35668) := x"10a0";
    tmp(35669) := x"10a0";
    tmp(35670) := x"1080";
    tmp(35671) := x"1080";
    tmp(35672) := x"1080";
    tmp(35673) := x"0880";
    tmp(35674) := x"0880";
    tmp(35675) := x"0860";
    tmp(35676) := x"0860";
    tmp(35677) := x"0860";
    tmp(35678) := x"0860";
    tmp(35679) := x"0860";
    tmp(35680) := x"1060";
    tmp(35681) := x"1060";
    tmp(35682) := x"1060";
    tmp(35683) := x"1060";
    tmp(35684) := x"1060";
    tmp(35685) := x"1060";
    tmp(35686) := x"1060";
    tmp(35687) := x"1040";
    tmp(35688) := x"1040";
    tmp(35689) := x"1040";
    tmp(35690) := x"1040";
    tmp(35691) := x"1040";
    tmp(35692) := x"0840";
    tmp(35693) := x"1040";
    tmp(35694) := x"1040";
    tmp(35695) := x"1040";
    tmp(35696) := x"1040";
    tmp(35697) := x"1040";
    tmp(35698) := x"1040";
    tmp(35699) := x"1040";
    tmp(35700) := x"1040";
    tmp(35701) := x"1040";
    tmp(35702) := x"1040";
    tmp(35703) := x"1040";
    tmp(35704) := x"1040";
    tmp(35705) := x"1040";
    tmp(35706) := x"1040";
    tmp(35707) := x"1040";
    tmp(35708) := x"1040";
    tmp(35709) := x"1040";
    tmp(35710) := x"1040";
    tmp(35711) := x"1040";
    tmp(35712) := x"0840";
    tmp(35713) := x"0840";
    tmp(35714) := x"1040";
    tmp(35715) := x"0840";
    tmp(35716) := x"0840";
    tmp(35717) := x"07e0";
    tmp(35718) := x"07e0";
    tmp(35719) := x"07e0";
    tmp(35720) := x"07e0";
    tmp(35721) := x"07e0";
    tmp(35722) := x"07e0";
    tmp(35723) := x"07e0";
    tmp(35724) := x"07e0";
    tmp(35725) := x"07e0";
    tmp(35726) := x"07e0";
    tmp(35727) := x"07e0";
    tmp(35728) := x"07e0";
    tmp(35729) := x"07e0";
    tmp(35730) := x"07e0";
    tmp(35731) := x"07e0";
    tmp(35732) := x"07e0";
    tmp(35733) := x"07e0";
    tmp(35734) := x"07e0";
    tmp(35735) := x"07e0";
    tmp(35736) := x"07e0";
    tmp(35737) := x"07e0";
    tmp(35738) := x"07e0";
    tmp(35739) := x"07e0";
    tmp(35740) := x"07e0";
    tmp(35741) := x"07e0";
    tmp(35742) := x"07e0";
    tmp(35743) := x"07e0";
    tmp(35744) := x"07e0";
    tmp(35745) := x"07e0";
    tmp(35746) := x"07e0";
    tmp(35747) := x"07e0";
    tmp(35748) := x"07e0";
    tmp(35749) := x"07e0";
    tmp(35750) := x"07e0";
    tmp(35751) := x"07e0";
    tmp(35752) := x"07e0";
    tmp(35753) := x"07e0";
    tmp(35754) := x"07e0";
    tmp(35755) := x"07e0";
    tmp(35756) := x"07e0";
    tmp(35757) := x"0840";
    tmp(35758) := x"0840";
    tmp(35759) := x"0840";
    tmp(35760) := x"0020";
    tmp(35761) := x"00e5";
    tmp(35762) := x"00c4";
    tmp(35763) := x"0083";
    tmp(35764) := x"00c4";
    tmp(35765) := x"00e4";
    tmp(35766) := x"00c4";
    tmp(35767) := x"00a4";
    tmp(35768) := x"00c4";
    tmp(35769) := x"00c4";
    tmp(35770) := x"00e5";
    tmp(35771) := x"00e5";
    tmp(35772) := x"00e5";
    tmp(35773) := x"08e5";
    tmp(35774) := x"08e5";
    tmp(35775) := x"08e4";
    tmp(35776) := x"00c4";
    tmp(35777) := x"00a3";
    tmp(35778) := x"08e4";
    tmp(35779) := x"0926";
    tmp(35780) := x"0926";
    tmp(35781) := x"0905";
    tmp(35782) := x"0947";
    tmp(35783) := x"09a8";
    tmp(35784) := x"09c9";
    tmp(35785) := x"09c9";
    tmp(35786) := x"09c8";
    tmp(35787) := x"09c8";
    tmp(35788) := x"09c8";
    tmp(35789) := x"0987";
    tmp(35790) := x"0905";
    tmp(35791) := x"00a3";
    tmp(35792) := x"0061";
    tmp(35793) := x"0082";
    tmp(35794) := x"0925";
    tmp(35795) := x"0967";
    tmp(35796) := x"0987";
    tmp(35797) := x"09a7";
    tmp(35798) := x"1186";
    tmp(35799) := x"08c2";
    tmp(35800) := x"08a1";
    tmp(35801) := x"1121";
    tmp(35802) := x"1981";
    tmp(35803) := x"1161";
    tmp(35804) := x"1181";
    tmp(35805) := x"1161";
    tmp(35806) := x"1140";
    tmp(35807) := x"1140";
    tmp(35808) := x"1140";
    tmp(35809) := x"1120";
    tmp(35810) := x"1140";
    tmp(35811) := x"1120";
    tmp(35812) := x"1120";
    tmp(35813) := x"0920";
    tmp(35814) := x"0940";
    tmp(35815) := x"1140";
    tmp(35816) := x"1140";
    tmp(35817) := x"1120";
    tmp(35818) := x"1140";
    tmp(35819) := x"1120";
    tmp(35820) := x"1140";
    tmp(35821) := x"1140";
    tmp(35822) := x"1120";
    tmp(35823) := x"1120";
    tmp(35824) := x"1120";
    tmp(35825) := x"0920";
    tmp(35826) := x"0920";
    tmp(35827) := x"0920";
    tmp(35828) := x"0920";
    tmp(35829) := x"0920";
    tmp(35830) := x"0920";
    tmp(35831) := x"0920";
    tmp(35832) := x"0920";
    tmp(35833) := x"0920";
    tmp(35834) := x"0900";
    tmp(35835) := x"0900";
    tmp(35836) := x"0900";
    tmp(35837) := x"0900";
    tmp(35838) := x"0900";
    tmp(35839) := x"0900";
    tmp(35840) := x"1101";
    tmp(35841) := x"1101";
    tmp(35842) := x"1121";
    tmp(35843) := x"1121";
    tmp(35844) := x"1121";
    tmp(35845) := x"1121";
    tmp(35846) := x"1121";
    tmp(35847) := x"1122";
    tmp(35848) := x"1102";
    tmp(35849) := x"1102";
    tmp(35850) := x"1102";
    tmp(35851) := x"1102";
    tmp(35852) := x"1102";
    tmp(35853) := x"1902";
    tmp(35854) := x"1901";
    tmp(35855) := x"1921";
    tmp(35856) := x"1921";
    tmp(35857) := x"1921";
    tmp(35858) := x"1921";
    tmp(35859) := x"1921";
    tmp(35860) := x"1941";
    tmp(35861) := x"1921";
    tmp(35862) := x"1941";
    tmp(35863) := x"1121";
    tmp(35864) := x"1121";
    tmp(35865) := x"1101";
    tmp(35866) := x"1101";
    tmp(35867) := x"0900";
    tmp(35868) := x"08e0";
    tmp(35869) := x"08e0";
    tmp(35870) := x"08e0";
    tmp(35871) := x"1100";
    tmp(35872) := x"0900";
    tmp(35873) := x"1100";
    tmp(35874) := x"1100";
    tmp(35875) := x"10e0";
    tmp(35876) := x"10e0";
    tmp(35877) := x"1100";
    tmp(35878) := x"1100";
    tmp(35879) := x"1101";
    tmp(35880) := x"1101";
    tmp(35881) := x"10e1";
    tmp(35882) := x"10e0";
    tmp(35883) := x"1100";
    tmp(35884) := x"1100";
    tmp(35885) := x"10e0";
    tmp(35886) := x"1100";
    tmp(35887) := x"1120";
    tmp(35888) := x"1120";
    tmp(35889) := x"1120";
    tmp(35890) := x"1120";
    tmp(35891) := x"0900";
    tmp(35892) := x"0900";
    tmp(35893) := x"0900";
    tmp(35894) := x"0920";
    tmp(35895) := x"0900";
    tmp(35896) := x"0900";
    tmp(35897) := x"0900";
    tmp(35898) := x"08e0";
    tmp(35899) := x"08e0";
    tmp(35900) := x"08e0";
    tmp(35901) := x"08c0";
    tmp(35902) := x"08c0";
    tmp(35903) := x"08c0";
    tmp(35904) := x"08c0";
    tmp(35905) := x"08a0";
    tmp(35906) := x"08a0";
    tmp(35907) := x"10a0";
    tmp(35908) := x"10a0";
    tmp(35909) := x"10a0";
    tmp(35910) := x"1080";
    tmp(35911) := x"1080";
    tmp(35912) := x"0880";
    tmp(35913) := x"0880";
    tmp(35914) := x"0880";
    tmp(35915) := x"0860";
    tmp(35916) := x"0860";
    tmp(35917) := x"0860";
    tmp(35918) := x"0860";
    tmp(35919) := x"0860";
    tmp(35920) := x"1060";
    tmp(35921) := x"1060";
    tmp(35922) := x"1060";
    tmp(35923) := x"1060";
    tmp(35924) := x"1040";
    tmp(35925) := x"1060";
    tmp(35926) := x"1060";
    tmp(35927) := x"1040";
    tmp(35928) := x"1040";
    tmp(35929) := x"1040";
    tmp(35930) := x"1040";
    tmp(35931) := x"0840";
    tmp(35932) := x"0840";
    tmp(35933) := x"1040";
    tmp(35934) := x"1040";
    tmp(35935) := x"1040";
    tmp(35936) := x"1040";
    tmp(35937) := x"1040";
    tmp(35938) := x"1040";
    tmp(35939) := x"1040";
    tmp(35940) := x"1040";
    tmp(35941) := x"1040";
    tmp(35942) := x"1040";
    tmp(35943) := x"1040";
    tmp(35944) := x"1040";
    tmp(35945) := x"1040";
    tmp(35946) := x"1040";
    tmp(35947) := x"1040";
    tmp(35948) := x"1040";
    tmp(35949) := x"1040";
    tmp(35950) := x"0840";
    tmp(35951) := x"1040";
    tmp(35952) := x"1040";
    tmp(35953) := x"1040";
    tmp(35954) := x"1040";
    tmp(35955) := x"1040";
    tmp(35956) := x"0840";
    tmp(35957) := x"07e0";
    tmp(35958) := x"07e0";
    tmp(35959) := x"07e0";
    tmp(35960) := x"07e0";
    tmp(35961) := x"07e0";
    tmp(35962) := x"07e0";
    tmp(35963) := x"07e0";
    tmp(35964) := x"07e0";
    tmp(35965) := x"07e0";
    tmp(35966) := x"07e0";
    tmp(35967) := x"07e0";
    tmp(35968) := x"07e0";
    tmp(35969) := x"07e0";
    tmp(35970) := x"07e0";
    tmp(35971) := x"07e0";
    tmp(35972) := x"07e0";
    tmp(35973) := x"07e0";
    tmp(35974) := x"07e0";
    tmp(35975) := x"07e0";
    tmp(35976) := x"07e0";
    tmp(35977) := x"07e0";
    tmp(35978) := x"07e0";
    tmp(35979) := x"07e0";
    tmp(35980) := x"07e0";
    tmp(35981) := x"07e0";
    tmp(35982) := x"07e0";
    tmp(35983) := x"07e0";
    tmp(35984) := x"07e0";
    tmp(35985) := x"07e0";
    tmp(35986) := x"07e0";
    tmp(35987) := x"07e0";
    tmp(35988) := x"07e0";
    tmp(35989) := x"07e0";
    tmp(35990) := x"07e0";
    tmp(35991) := x"07e0";
    tmp(35992) := x"07e0";
    tmp(35993) := x"07e0";
    tmp(35994) := x"07e0";
    tmp(35995) := x"07e0";
    tmp(35996) := x"07e0";
    tmp(35997) := x"0840";
    tmp(35998) := x"0840";
    tmp(35999) := x"0840";
    tmp(36000) := x"0020";
    tmp(36001) := x"00c4";
    tmp(36002) := x"00a3";
    tmp(36003) := x"00a3";
    tmp(36004) := x"00c4";
    tmp(36005) := x"0905";
    tmp(36006) := x"00e4";
    tmp(36007) := x"00c4";
    tmp(36008) := x"00a3";
    tmp(36009) := x"00a3";
    tmp(36010) := x"00a3";
    tmp(36011) := x"00c4";
    tmp(36012) := x"00c4";
    tmp(36013) := x"00c4";
    tmp(36014) := x"08e5";
    tmp(36015) := x"08e5";
    tmp(36016) := x"08e5";
    tmp(36017) := x"08e5";
    tmp(36018) := x"08c4";
    tmp(36019) := x"08a3";
    tmp(36020) := x"00a3";
    tmp(36021) := x"08e4";
    tmp(36022) := x"0987";
    tmp(36023) := x"09a8";
    tmp(36024) := x"09a8";
    tmp(36025) := x"0987";
    tmp(36026) := x"0987";
    tmp(36027) := x"0967";
    tmp(36028) := x"0905";
    tmp(36029) := x"00c3";
    tmp(36030) := x"00a2";
    tmp(36031) := x"00e3";
    tmp(36032) := x"09c7";
    tmp(36033) := x"11e9";
    tmp(36034) := x"0925";
    tmp(36035) := x"08e4";
    tmp(36036) := x"08e3";
    tmp(36037) := x"08c2";
    tmp(36038) := x"0061";
    tmp(36039) := x"08c1";
    tmp(36040) := x"1161";
    tmp(36041) := x"1181";
    tmp(36042) := x"1161";
    tmp(36043) := x"1161";
    tmp(36044) := x"1161";
    tmp(36045) := x"1161";
    tmp(36046) := x"1140";
    tmp(36047) := x"1120";
    tmp(36048) := x"1120";
    tmp(36049) := x"1120";
    tmp(36050) := x"1120";
    tmp(36051) := x"0920";
    tmp(36052) := x"1140";
    tmp(36053) := x"1120";
    tmp(36054) := x"1140";
    tmp(36055) := x"0940";
    tmp(36056) := x"0920";
    tmp(36057) := x"1120";
    tmp(36058) := x"1120";
    tmp(36059) := x"1140";
    tmp(36060) := x"1140";
    tmp(36061) := x"0920";
    tmp(36062) := x"1120";
    tmp(36063) := x"1120";
    tmp(36064) := x"1120";
    tmp(36065) := x"1120";
    tmp(36066) := x"0920";
    tmp(36067) := x"1120";
    tmp(36068) := x"1120";
    tmp(36069) := x"1120";
    tmp(36070) := x"0920";
    tmp(36071) := x"0920";
    tmp(36072) := x"0920";
    tmp(36073) := x"0920";
    tmp(36074) := x"0920";
    tmp(36075) := x"0900";
    tmp(36076) := x"0900";
    tmp(36077) := x"0900";
    tmp(36078) := x"0900";
    tmp(36079) := x"0900";
    tmp(36080) := x"0920";
    tmp(36081) := x"1121";
    tmp(36082) := x"1121";
    tmp(36083) := x"1121";
    tmp(36084) := x"1121";
    tmp(36085) := x"1121";
    tmp(36086) := x"1101";
    tmp(36087) := x"1121";
    tmp(36088) := x"1121";
    tmp(36089) := x"1102";
    tmp(36090) := x"1101";
    tmp(36091) := x"1101";
    tmp(36092) := x"1101";
    tmp(36093) := x"1101";
    tmp(36094) := x"1901";
    tmp(36095) := x"1921";
    tmp(36096) := x"1921";
    tmp(36097) := x"1921";
    tmp(36098) := x"1921";
    tmp(36099) := x"1941";
    tmp(36100) := x"1941";
    tmp(36101) := x"1941";
    tmp(36102) := x"1121";
    tmp(36103) := x"1121";
    tmp(36104) := x"1101";
    tmp(36105) := x"1121";
    tmp(36106) := x"0900";
    tmp(36107) := x"0900";
    tmp(36108) := x"08e0";
    tmp(36109) := x"08e0";
    tmp(36110) := x"08e0";
    tmp(36111) := x"0900";
    tmp(36112) := x"0900";
    tmp(36113) := x"1100";
    tmp(36114) := x"0900";
    tmp(36115) := x"08e0";
    tmp(36116) := x"10e0";
    tmp(36117) := x"1100";
    tmp(36118) := x"1100";
    tmp(36119) := x"1101";
    tmp(36120) := x"1101";
    tmp(36121) := x"10e1";
    tmp(36122) := x"10e1";
    tmp(36123) := x"1100";
    tmp(36124) := x"10e0";
    tmp(36125) := x"08e0";
    tmp(36126) := x"1100";
    tmp(36127) := x"1120";
    tmp(36128) := x"1120";
    tmp(36129) := x"1120";
    tmp(36130) := x"0920";
    tmp(36131) := x"0900";
    tmp(36132) := x"0900";
    tmp(36133) := x"0920";
    tmp(36134) := x"0920";
    tmp(36135) := x"0920";
    tmp(36136) := x"0900";
    tmp(36137) := x"0900";
    tmp(36138) := x"08e0";
    tmp(36139) := x"08e0";
    tmp(36140) := x"08e0";
    tmp(36141) := x"08c0";
    tmp(36142) := x"08c0";
    tmp(36143) := x"08c0";
    tmp(36144) := x"08c0";
    tmp(36145) := x"08a0";
    tmp(36146) := x"08a0";
    tmp(36147) := x"08a0";
    tmp(36148) := x"10a0";
    tmp(36149) := x"10a0";
    tmp(36150) := x"1080";
    tmp(36151) := x"0880";
    tmp(36152) := x"0880";
    tmp(36153) := x"0880";
    tmp(36154) := x"0880";
    tmp(36155) := x"0880";
    tmp(36156) := x"0860";
    tmp(36157) := x"0860";
    tmp(36158) := x"0860";
    tmp(36159) := x"0860";
    tmp(36160) := x"1060";
    tmp(36161) := x"1060";
    tmp(36162) := x"1060";
    tmp(36163) := x"1060";
    tmp(36164) := x"1060";
    tmp(36165) := x"1060";
    tmp(36166) := x"1060";
    tmp(36167) := x"1040";
    tmp(36168) := x"1040";
    tmp(36169) := x"1040";
    tmp(36170) := x"1040";
    tmp(36171) := x"1040";
    tmp(36172) := x"1040";
    tmp(36173) := x"1040";
    tmp(36174) := x"1040";
    tmp(36175) := x"1040";
    tmp(36176) := x"1040";
    tmp(36177) := x"1040";
    tmp(36178) := x"1040";
    tmp(36179) := x"1040";
    tmp(36180) := x"1040";
    tmp(36181) := x"1040";
    tmp(36182) := x"1060";
    tmp(36183) := x"1040";
    tmp(36184) := x"1040";
    tmp(36185) := x"1040";
    tmp(36186) := x"1040";
    tmp(36187) := x"1040";
    tmp(36188) := x"1040";
    tmp(36189) := x"1040";
    tmp(36190) := x"1040";
    tmp(36191) := x"1040";
    tmp(36192) := x"1040";
    tmp(36193) := x"1040";
    tmp(36194) := x"0840";
    tmp(36195) := x"1040";
    tmp(36196) := x"0840";
    tmp(36197) := x"07e0";
    tmp(36198) := x"07e0";
    tmp(36199) := x"07e0";
    tmp(36200) := x"07e0";
    tmp(36201) := x"07e0";
    tmp(36202) := x"07e0";
    tmp(36203) := x"07e0";
    tmp(36204) := x"07e0";
    tmp(36205) := x"07e0";
    tmp(36206) := x"07e0";
    tmp(36207) := x"07e0";
    tmp(36208) := x"07e0";
    tmp(36209) := x"07e0";
    tmp(36210) := x"07e0";
    tmp(36211) := x"07e0";
    tmp(36212) := x"07e0";
    tmp(36213) := x"07e0";
    tmp(36214) := x"07e0";
    tmp(36215) := x"07e0";
    tmp(36216) := x"07e0";
    tmp(36217) := x"07e0";
    tmp(36218) := x"07e0";
    tmp(36219) := x"07e0";
    tmp(36220) := x"07e0";
    tmp(36221) := x"07e0";
    tmp(36222) := x"07e0";
    tmp(36223) := x"07e0";
    tmp(36224) := x"07e0";
    tmp(36225) := x"07e0";
    tmp(36226) := x"07e0";
    tmp(36227) := x"07e0";
    tmp(36228) := x"07e0";
    tmp(36229) := x"07e0";
    tmp(36230) := x"07e0";
    tmp(36231) := x"07e0";
    tmp(36232) := x"07e0";
    tmp(36233) := x"07e0";
    tmp(36234) := x"07e0";
    tmp(36235) := x"07e0";
    tmp(36236) := x"07e0";
    tmp(36237) := x"0840";
    tmp(36238) := x"0840";
    tmp(36239) := x"0840";
    tmp(36240) := x"0020";
    tmp(36241) := x"00c4";
    tmp(36242) := x"00a3";
    tmp(36243) := x"0082";
    tmp(36244) := x"0082";
    tmp(36245) := x"00c4";
    tmp(36246) := x"08e5";
    tmp(36247) := x"08e5";
    tmp(36248) := x"00c4";
    tmp(36249) := x"00c4";
    tmp(36250) := x"00c4";
    tmp(36251) := x"00c3";
    tmp(36252) := x"00c3";
    tmp(36253) := x"00a3";
    tmp(36254) := x"00a3";
    tmp(36255) := x"00a3";
    tmp(36256) := x"00a3";
    tmp(36257) := x"00a4";
    tmp(36258) := x"00a4";
    tmp(36259) := x"00c4";
    tmp(36260) := x"0905";
    tmp(36261) := x"0946";
    tmp(36262) := x"0967";
    tmp(36263) := x"09a8";
    tmp(36264) := x"09a8";
    tmp(36265) := x"0967";
    tmp(36266) := x"0946";
    tmp(36267) := x"0925";
    tmp(36268) := x"00e4";
    tmp(36269) := x"0925";
    tmp(36270) := x"0a09";
    tmp(36271) := x"124a";
    tmp(36272) := x"09a7";
    tmp(36273) := x"08c3";
    tmp(36274) := x"0041";
    tmp(36275) := x"0020";
    tmp(36276) := x"0040";
    tmp(36277) := x"0860";
    tmp(36278) := x"0901";
    tmp(36279) := x"1181";
    tmp(36280) := x"1181";
    tmp(36281) := x"1181";
    tmp(36282) := x"1161";
    tmp(36283) := x"1161";
    tmp(36284) := x"1161";
    tmp(36285) := x"1161";
    tmp(36286) := x"1140";
    tmp(36287) := x"1120";
    tmp(36288) := x"0920";
    tmp(36289) := x"0920";
    tmp(36290) := x"0920";
    tmp(36291) := x"0920";
    tmp(36292) := x"0920";
    tmp(36293) := x"1120";
    tmp(36294) := x"1120";
    tmp(36295) := x"0920";
    tmp(36296) := x"1140";
    tmp(36297) := x"1120";
    tmp(36298) := x"1140";
    tmp(36299) := x"1140";
    tmp(36300) := x"1140";
    tmp(36301) := x"1120";
    tmp(36302) := x"1120";
    tmp(36303) := x"1140";
    tmp(36304) := x"1120";
    tmp(36305) := x"1120";
    tmp(36306) := x"1120";
    tmp(36307) := x"1120";
    tmp(36308) := x"1120";
    tmp(36309) := x"1120";
    tmp(36310) := x"1120";
    tmp(36311) := x"1120";
    tmp(36312) := x"0920";
    tmp(36313) := x"0920";
    tmp(36314) := x"0920";
    tmp(36315) := x"0920";
    tmp(36316) := x"0900";
    tmp(36317) := x"0900";
    tmp(36318) := x"0900";
    tmp(36319) := x"0900";
    tmp(36320) := x"0900";
    tmp(36321) := x"1121";
    tmp(36322) := x"1121";
    tmp(36323) := x"1121";
    tmp(36324) := x"1121";
    tmp(36325) := x"1121";
    tmp(36326) := x"1121";
    tmp(36327) := x"1121";
    tmp(36328) := x"1121";
    tmp(36329) := x"1101";
    tmp(36330) := x"1101";
    tmp(36331) := x"1101";
    tmp(36332) := x"1101";
    tmp(36333) := x"1101";
    tmp(36334) := x"1121";
    tmp(36335) := x"1921";
    tmp(36336) := x"1921";
    tmp(36337) := x"1921";
    tmp(36338) := x"1941";
    tmp(36339) := x"1941";
    tmp(36340) := x"1941";
    tmp(36341) := x"1941";
    tmp(36342) := x"1121";
    tmp(36343) := x"1121";
    tmp(36344) := x"1101";
    tmp(36345) := x"1101";
    tmp(36346) := x"08e0";
    tmp(36347) := x"08e0";
    tmp(36348) := x"08e0";
    tmp(36349) := x"08e0";
    tmp(36350) := x"08e0";
    tmp(36351) := x"0900";
    tmp(36352) := x"0900";
    tmp(36353) := x"0900";
    tmp(36354) := x"08e0";
    tmp(36355) := x"08e0";
    tmp(36356) := x"10e0";
    tmp(36357) := x"10e0";
    tmp(36358) := x"1100";
    tmp(36359) := x"1101";
    tmp(36360) := x"10e0";
    tmp(36361) := x"10e0";
    tmp(36362) := x"10e0";
    tmp(36363) := x"08e0";
    tmp(36364) := x"08e0";
    tmp(36365) := x"08e0";
    tmp(36366) := x"08e0";
    tmp(36367) := x"1100";
    tmp(36368) := x"1120";
    tmp(36369) := x"1120";
    tmp(36370) := x"0920";
    tmp(36371) := x"0900";
    tmp(36372) := x"0900";
    tmp(36373) := x"0920";
    tmp(36374) := x"0920";
    tmp(36375) := x"0900";
    tmp(36376) := x"0900";
    tmp(36377) := x"0900";
    tmp(36378) := x"08e0";
    tmp(36379) := x"08e0";
    tmp(36380) := x"08e0";
    tmp(36381) := x"08c0";
    tmp(36382) := x"08c0";
    tmp(36383) := x"08c0";
    tmp(36384) := x"08a0";
    tmp(36385) := x"08a0";
    tmp(36386) := x"08a0";
    tmp(36387) := x"08a0";
    tmp(36388) := x"10a0";
    tmp(36389) := x"0880";
    tmp(36390) := x"0880";
    tmp(36391) := x"0880";
    tmp(36392) := x"0880";
    tmp(36393) := x"0880";
    tmp(36394) := x"0880";
    tmp(36395) := x"0880";
    tmp(36396) := x"0860";
    tmp(36397) := x"0860";
    tmp(36398) := x"1060";
    tmp(36399) := x"1060";
    tmp(36400) := x"1060";
    tmp(36401) := x"1060";
    tmp(36402) := x"1060";
    tmp(36403) := x"1060";
    tmp(36404) := x"1060";
    tmp(36405) := x"1060";
    tmp(36406) := x"1060";
    tmp(36407) := x"1060";
    tmp(36408) := x"1040";
    tmp(36409) := x"1040";
    tmp(36410) := x"1040";
    tmp(36411) := x"1040";
    tmp(36412) := x"1040";
    tmp(36413) := x"1040";
    tmp(36414) := x"1040";
    tmp(36415) := x"1040";
    tmp(36416) := x"1040";
    tmp(36417) := x"1040";
    tmp(36418) := x"1040";
    tmp(36419) := x"1040";
    tmp(36420) := x"1060";
    tmp(36421) := x"1060";
    tmp(36422) := x"1040";
    tmp(36423) := x"1060";
    tmp(36424) := x"1060";
    tmp(36425) := x"1060";
    tmp(36426) := x"1060";
    tmp(36427) := x"1040";
    tmp(36428) := x"1040";
    tmp(36429) := x"1040";
    tmp(36430) := x"1040";
    tmp(36431) := x"1040";
    tmp(36432) := x"1040";
    tmp(36433) := x"0840";
    tmp(36434) := x"1040";
    tmp(36435) := x"1040";
    tmp(36436) := x"1040";
    tmp(36437) := x"07e0";
    tmp(36438) := x"07e0";
    tmp(36439) := x"07e0";
    tmp(36440) := x"07e0";
    tmp(36441) := x"07e0";
    tmp(36442) := x"07e0";
    tmp(36443) := x"07e0";
    tmp(36444) := x"07e0";
    tmp(36445) := x"07e0";
    tmp(36446) := x"07e0";
    tmp(36447) := x"07e0";
    tmp(36448) := x"07e0";
    tmp(36449) := x"07e0";
    tmp(36450) := x"07e0";
    tmp(36451) := x"07e0";
    tmp(36452) := x"07e0";
    tmp(36453) := x"07e0";
    tmp(36454) := x"07e0";
    tmp(36455) := x"07e0";
    tmp(36456) := x"07e0";
    tmp(36457) := x"07e0";
    tmp(36458) := x"07e0";
    tmp(36459) := x"07e0";
    tmp(36460) := x"07e0";
    tmp(36461) := x"07e0";
    tmp(36462) := x"07e0";
    tmp(36463) := x"07e0";
    tmp(36464) := x"07e0";
    tmp(36465) := x"07e0";
    tmp(36466) := x"07e0";
    tmp(36467) := x"07e0";
    tmp(36468) := x"07e0";
    tmp(36469) := x"07e0";
    tmp(36470) := x"07e0";
    tmp(36471) := x"07e0";
    tmp(36472) := x"07e0";
    tmp(36473) := x"07e0";
    tmp(36474) := x"07e0";
    tmp(36475) := x"07e0";
    tmp(36476) := x"07e0";
    tmp(36477) := x"0840";
    tmp(36478) := x"0840";
    tmp(36479) := x"0840";
    tmp(36480) := x"0020";
    tmp(36481) := x"00e5";
    tmp(36482) := x"00c4";
    tmp(36483) := x"00c3";
    tmp(36484) := x"0083";
    tmp(36485) := x"0083";
    tmp(36486) := x"00c3";
    tmp(36487) := x"00e4";
    tmp(36488) := x"0925";
    tmp(36489) := x"0925";
    tmp(36490) := x"0905";
    tmp(36491) := x"08e5";
    tmp(36492) := x"08e5";
    tmp(36493) := x"08e5";
    tmp(36494) := x"0905";
    tmp(36495) := x"0905";
    tmp(36496) := x"0926";
    tmp(36497) := x"0947";
    tmp(36498) := x"09a8";
    tmp(36499) := x"09c9";
    tmp(36500) := x"09ea";
    tmp(36501) := x"09c9";
    tmp(36502) := x"0966";
    tmp(36503) := x"0925";
    tmp(36504) := x"0904";
    tmp(36505) := x"0925";
    tmp(36506) := x"0925";
    tmp(36507) := x"0905";
    tmp(36508) := x"09a8";
    tmp(36509) := x"0a2b";
    tmp(36510) := x"09c9";
    tmp(36511) := x"08a3";
    tmp(36512) := x"0041";
    tmp(36513) := x"0020";
    tmp(36514) := x"0020";
    tmp(36515) := x"0020";
    tmp(36516) := x"0880";
    tmp(36517) := x"1121";
    tmp(36518) := x"1161";
    tmp(36519) := x"1161";
    tmp(36520) := x"1161";
    tmp(36521) := x"1161";
    tmp(36522) := x"1161";
    tmp(36523) := x"1141";
    tmp(36524) := x"1161";
    tmp(36525) := x"1140";
    tmp(36526) := x"1140";
    tmp(36527) := x"1140";
    tmp(36528) := x"1120";
    tmp(36529) := x"1120";
    tmp(36530) := x"1120";
    tmp(36531) := x"0920";
    tmp(36532) := x"1120";
    tmp(36533) := x"1120";
    tmp(36534) := x"1120";
    tmp(36535) := x"1140";
    tmp(36536) := x"1140";
    tmp(36537) := x"1140";
    tmp(36538) := x"1120";
    tmp(36539) := x"1140";
    tmp(36540) := x"1140";
    tmp(36541) := x"1120";
    tmp(36542) := x"1120";
    tmp(36543) := x"1140";
    tmp(36544) := x"1140";
    tmp(36545) := x"1120";
    tmp(36546) := x"1140";
    tmp(36547) := x"1140";
    tmp(36548) := x"1140";
    tmp(36549) := x"1120";
    tmp(36550) := x"1120";
    tmp(36551) := x"1120";
    tmp(36552) := x"1120";
    tmp(36553) := x"0920";
    tmp(36554) := x"0920";
    tmp(36555) := x"0920";
    tmp(36556) := x"0920";
    tmp(36557) := x"0900";
    tmp(36558) := x"0900";
    tmp(36559) := x"0900";
    tmp(36560) := x"0900";
    tmp(36561) := x"0900";
    tmp(36562) := x"0900";
    tmp(36563) := x"1101";
    tmp(36564) := x"1121";
    tmp(36565) := x"1121";
    tmp(36566) := x"1101";
    tmp(36567) := x"1121";
    tmp(36568) := x"1121";
    tmp(36569) := x"1101";
    tmp(36570) := x"1101";
    tmp(36571) := x"1101";
    tmp(36572) := x"1101";
    tmp(36573) := x"1101";
    tmp(36574) := x"1921";
    tmp(36575) := x"1121";
    tmp(36576) := x"1921";
    tmp(36577) := x"1941";
    tmp(36578) := x"1941";
    tmp(36579) := x"1941";
    tmp(36580) := x"1141";
    tmp(36581) := x"1141";
    tmp(36582) := x"1121";
    tmp(36583) := x"1121";
    tmp(36584) := x"1121";
    tmp(36585) := x"0900";
    tmp(36586) := x"0900";
    tmp(36587) := x"08e0";
    tmp(36588) := x"08e0";
    tmp(36589) := x"0900";
    tmp(36590) := x"08e0";
    tmp(36591) := x"08e0";
    tmp(36592) := x"0900";
    tmp(36593) := x"08e0";
    tmp(36594) := x"08e0";
    tmp(36595) := x"08e0";
    tmp(36596) := x"08e0";
    tmp(36597) := x"10e0";
    tmp(36598) := x"1100";
    tmp(36599) := x"1100";
    tmp(36600) := x"10e0";
    tmp(36601) := x"1101";
    tmp(36602) := x"10e0";
    tmp(36603) := x"08c0";
    tmp(36604) := x"08e0";
    tmp(36605) := x"08e0";
    tmp(36606) := x"08e0";
    tmp(36607) := x"1100";
    tmp(36608) := x"1100";
    tmp(36609) := x"1120";
    tmp(36610) := x"0920";
    tmp(36611) := x"0900";
    tmp(36612) := x"0900";
    tmp(36613) := x"0900";
    tmp(36614) := x"0920";
    tmp(36615) := x"0920";
    tmp(36616) := x"0900";
    tmp(36617) := x"0900";
    tmp(36618) := x"0900";
    tmp(36619) := x"08e0";
    tmp(36620) := x"08e0";
    tmp(36621) := x"08c0";
    tmp(36622) := x"08c0";
    tmp(36623) := x"08c0";
    tmp(36624) := x"08c0";
    tmp(36625) := x"08a0";
    tmp(36626) := x"08a0";
    tmp(36627) := x"08a0";
    tmp(36628) := x"08a0";
    tmp(36629) := x"0880";
    tmp(36630) := x"0880";
    tmp(36631) := x"0880";
    tmp(36632) := x"0880";
    tmp(36633) := x"0880";
    tmp(36634) := x"0880";
    tmp(36635) := x"0880";
    tmp(36636) := x"1060";
    tmp(36637) := x"1060";
    tmp(36638) := x"1060";
    tmp(36639) := x"1060";
    tmp(36640) := x"1060";
    tmp(36641) := x"1060";
    tmp(36642) := x"1060";
    tmp(36643) := x"1060";
    tmp(36644) := x"1060";
    tmp(36645) := x"1060";
    tmp(36646) := x"1060";
    tmp(36647) := x"1060";
    tmp(36648) := x"1040";
    tmp(36649) := x"1040";
    tmp(36650) := x"1040";
    tmp(36651) := x"1040";
    tmp(36652) := x"1040";
    tmp(36653) := x"1040";
    tmp(36654) := x"1040";
    tmp(36655) := x"1040";
    tmp(36656) := x"1040";
    tmp(36657) := x"1060";
    tmp(36658) := x"1060";
    tmp(36659) := x"1040";
    tmp(36660) := x"1040";
    tmp(36661) := x"1040";
    tmp(36662) := x"1040";
    tmp(36663) := x"1060";
    tmp(36664) := x"1060";
    tmp(36665) := x"1060";
    tmp(36666) := x"1060";
    tmp(36667) := x"1060";
    tmp(36668) := x"1060";
    tmp(36669) := x"1060";
    tmp(36670) := x"1040";
    tmp(36671) := x"1040";
    tmp(36672) := x"1060";
    tmp(36673) := x"1040";
    tmp(36674) := x"1040";
    tmp(36675) := x"1040";
    tmp(36676) := x"0840";
    tmp(36677) := x"07e0";
    tmp(36678) := x"07e0";
    tmp(36679) := x"07e0";
    tmp(36680) := x"07e0";
    tmp(36681) := x"07e0";
    tmp(36682) := x"07e0";
    tmp(36683) := x"07e0";
    tmp(36684) := x"07e0";
    tmp(36685) := x"07e0";
    tmp(36686) := x"07e0";
    tmp(36687) := x"07e0";
    tmp(36688) := x"07e0";
    tmp(36689) := x"07e0";
    tmp(36690) := x"07e0";
    tmp(36691) := x"07e0";
    tmp(36692) := x"07e0";
    tmp(36693) := x"07e0";
    tmp(36694) := x"07e0";
    tmp(36695) := x"07e0";
    tmp(36696) := x"07e0";
    tmp(36697) := x"07e0";
    tmp(36698) := x"07e0";
    tmp(36699) := x"07e0";
    tmp(36700) := x"07e0";
    tmp(36701) := x"07e0";
    tmp(36702) := x"07e0";
    tmp(36703) := x"07e0";
    tmp(36704) := x"07e0";
    tmp(36705) := x"07e0";
    tmp(36706) := x"07e0";
    tmp(36707) := x"07e0";
    tmp(36708) := x"07e0";
    tmp(36709) := x"07e0";
    tmp(36710) := x"07e0";
    tmp(36711) := x"07e0";
    tmp(36712) := x"07e0";
    tmp(36713) := x"07e0";
    tmp(36714) := x"07e0";
    tmp(36715) := x"07e0";
    tmp(36716) := x"07e0";
    tmp(36717) := x"0840";
    tmp(36718) := x"0840";
    tmp(36719) := x"0840";
    tmp(36720) := x"0020";
    tmp(36721) := x"0105";
    tmp(36722) := x"00e4";
    tmp(36723) := x"00e4";
    tmp(36724) := x"00e4";
    tmp(36725) := x"00c4";
    tmp(36726) := x"00c4";
    tmp(36727) := x"00e5";
    tmp(36728) := x"0925";
    tmp(36729) := x"0905";
    tmp(36730) := x"0946";
    tmp(36731) := x"0988";
    tmp(36732) := x"0988";
    tmp(36733) := x"0968";
    tmp(36734) := x"09ea";
    tmp(36735) := x"0a0a";
    tmp(36736) := x"0a0b";
    tmp(36737) := x"0a0b";
    tmp(36738) := x"09e9";
    tmp(36739) := x"09a8";
    tmp(36740) := x"0967";
    tmp(36741) := x"0966";
    tmp(36742) := x"0966";
    tmp(36743) := x"0946";
    tmp(36744) := x"0945";
    tmp(36745) := x"00c3";
    tmp(36746) := x"00a3";
    tmp(36747) := x"0946";
    tmp(36748) := x"0a0a";
    tmp(36749) := x"0925";
    tmp(36750) := x"0061";
    tmp(36751) := x"0020";
    tmp(36752) := x"0020";
    tmp(36753) := x"0040";
    tmp(36754) := x"0880";
    tmp(36755) := x"08e1";
    tmp(36756) := x"1141";
    tmp(36757) := x"1141";
    tmp(36758) := x"1161";
    tmp(36759) := x"1161";
    tmp(36760) := x"1141";
    tmp(36761) := x"1141";
    tmp(36762) := x"1161";
    tmp(36763) := x"1161";
    tmp(36764) := x"1161";
    tmp(36765) := x"1161";
    tmp(36766) := x"1161";
    tmp(36767) := x"1140";
    tmp(36768) := x"1140";
    tmp(36769) := x"1120";
    tmp(36770) := x"0920";
    tmp(36771) := x"1120";
    tmp(36772) := x"1140";
    tmp(36773) := x"1140";
    tmp(36774) := x"1140";
    tmp(36775) := x"1140";
    tmp(36776) := x"1140";
    tmp(36777) := x"1140";
    tmp(36778) := x"1140";
    tmp(36779) := x"1140";
    tmp(36780) := x"1140";
    tmp(36781) := x"1140";
    tmp(36782) := x"1140";
    tmp(36783) := x"1140";
    tmp(36784) := x"1140";
    tmp(36785) := x"1140";
    tmp(36786) := x"1140";
    tmp(36787) := x"1140";
    tmp(36788) := x"1140";
    tmp(36789) := x"1140";
    tmp(36790) := x"1140";
    tmp(36791) := x"1120";
    tmp(36792) := x"1140";
    tmp(36793) := x"1120";
    tmp(36794) := x"0920";
    tmp(36795) := x"0920";
    tmp(36796) := x"0900";
    tmp(36797) := x"0920";
    tmp(36798) := x"0900";
    tmp(36799) := x"0900";
    tmp(36800) := x"0900";
    tmp(36801) := x"0900";
    tmp(36802) := x"0900";
    tmp(36803) := x"1121";
    tmp(36804) := x"1121";
    tmp(36805) := x"1121";
    tmp(36806) := x"1121";
    tmp(36807) := x"1121";
    tmp(36808) := x"1121";
    tmp(36809) := x"1101";
    tmp(36810) := x"1121";
    tmp(36811) := x"1101";
    tmp(36812) := x"1101";
    tmp(36813) := x"1121";
    tmp(36814) := x"1121";
    tmp(36815) := x"1121";
    tmp(36816) := x"1941";
    tmp(36817) := x"1941";
    tmp(36818) := x"1941";
    tmp(36819) := x"1141";
    tmp(36820) := x"1141";
    tmp(36821) := x"1121";
    tmp(36822) := x"1121";
    tmp(36823) := x"1121";
    tmp(36824) := x"0900";
    tmp(36825) := x"0900";
    tmp(36826) := x"0900";
    tmp(36827) := x"08e0";
    tmp(36828) := x"0900";
    tmp(36829) := x"08e0";
    tmp(36830) := x"08e0";
    tmp(36831) := x"08e0";
    tmp(36832) := x"08e0";
    tmp(36833) := x"08e0";
    tmp(36834) := x"08e0";
    tmp(36835) := x"08e0";
    tmp(36836) := x"08e0";
    tmp(36837) := x"10e0";
    tmp(36838) := x"1100";
    tmp(36839) := x"1100";
    tmp(36840) := x"1100";
    tmp(36841) := x"10e0";
    tmp(36842) := x"08c0";
    tmp(36843) := x"08c0";
    tmp(36844) := x"08c0";
    tmp(36845) := x"08e0";
    tmp(36846) := x"08e0";
    tmp(36847) := x"08e0";
    tmp(36848) := x"0900";
    tmp(36849) := x"0900";
    tmp(36850) := x"0900";
    tmp(36851) := x"0900";
    tmp(36852) := x"0900";
    tmp(36853) := x"0920";
    tmp(36854) := x"0920";
    tmp(36855) := x"0920";
    tmp(36856) := x"0900";
    tmp(36857) := x"0900";
    tmp(36858) := x"0900";
    tmp(36859) := x"08e0";
    tmp(36860) := x"08e0";
    tmp(36861) := x"08e0";
    tmp(36862) := x"08c0";
    tmp(36863) := x"08c0";
    tmp(36864) := x"08c0";
    tmp(36865) := x"08a0";
    tmp(36866) := x"08a0";
    tmp(36867) := x"08a0";
    tmp(36868) := x"08a0";
    tmp(36869) := x"0880";
    tmp(36870) := x"1080";
    tmp(36871) := x"0880";
    tmp(36872) := x"0880";
    tmp(36873) := x"0880";
    tmp(36874) := x"1080";
    tmp(36875) := x"1080";
    tmp(36876) := x"1080";
    tmp(36877) := x"1080";
    tmp(36878) := x"1080";
    tmp(36879) := x"1060";
    tmp(36880) := x"1060";
    tmp(36881) := x"1060";
    tmp(36882) := x"1060";
    tmp(36883) := x"1060";
    tmp(36884) := x"1060";
    tmp(36885) := x"1060";
    tmp(36886) := x"1060";
    tmp(36887) := x"1060";
    tmp(36888) := x"1060";
    tmp(36889) := x"1040";
    tmp(36890) := x"1040";
    tmp(36891) := x"1040";
    tmp(36892) := x"1040";
    tmp(36893) := x"1040";
    tmp(36894) := x"1040";
    tmp(36895) := x"1040";
    tmp(36896) := x"1040";
    tmp(36897) := x"1040";
    tmp(36898) := x"1060";
    tmp(36899) := x"1060";
    tmp(36900) := x"1060";
    tmp(36901) := x"1060";
    tmp(36902) := x"1060";
    tmp(36903) := x"1060";
    tmp(36904) := x"1060";
    tmp(36905) := x"1060";
    tmp(36906) := x"1060";
    tmp(36907) := x"1060";
    tmp(36908) := x"1060";
    tmp(36909) := x"1060";
    tmp(36910) := x"1060";
    tmp(36911) := x"1040";
    tmp(36912) := x"1040";
    tmp(36913) := x"1040";
    tmp(36914) := x"1040";
    tmp(36915) := x"1040";
    tmp(36916) := x"0840";
    tmp(36917) := x"07e0";
    tmp(36918) := x"07e0";
    tmp(36919) := x"07e0";
    tmp(36920) := x"07e0";
    tmp(36921) := x"07e0";
    tmp(36922) := x"07e0";
    tmp(36923) := x"07e0";
    tmp(36924) := x"07e0";
    tmp(36925) := x"07e0";
    tmp(36926) := x"07e0";
    tmp(36927) := x"07e0";
    tmp(36928) := x"07e0";
    tmp(36929) := x"07e0";
    tmp(36930) := x"07e0";
    tmp(36931) := x"07e0";
    tmp(36932) := x"07e0";
    tmp(36933) := x"07e0";
    tmp(36934) := x"07e0";
    tmp(36935) := x"07e0";
    tmp(36936) := x"07e0";
    tmp(36937) := x"07e0";
    tmp(36938) := x"07e0";
    tmp(36939) := x"07e0";
    tmp(36940) := x"07e0";
    tmp(36941) := x"07e0";
    tmp(36942) := x"07e0";
    tmp(36943) := x"07e0";
    tmp(36944) := x"07e0";
    tmp(36945) := x"07e0";
    tmp(36946) := x"07e0";
    tmp(36947) := x"07e0";
    tmp(36948) := x"07e0";
    tmp(36949) := x"07e0";
    tmp(36950) := x"07e0";
    tmp(36951) := x"07e0";
    tmp(36952) := x"07e0";
    tmp(36953) := x"07e0";
    tmp(36954) := x"07e0";
    tmp(36955) := x"07e0";
    tmp(36956) := x"07e0";
    tmp(36957) := x"0840";
    tmp(36958) := x"0840";
    tmp(36959) := x"0840";
    tmp(36960) := x"0020";
    tmp(36961) := x"00e4";
    tmp(36962) := x"0105";
    tmp(36963) := x"0925";
    tmp(36964) := x"0946";
    tmp(36965) := x"0946";
    tmp(36966) := x"0926";
    tmp(36967) := x"0926";
    tmp(36968) := x"0905";
    tmp(36969) := x"0926";
    tmp(36970) := x"0988";
    tmp(36971) := x"09ca";
    tmp(36972) := x"0988";
    tmp(36973) := x"0988";
    tmp(36974) := x"09ca";
    tmp(36975) := x"09a9";
    tmp(36976) := x"0988";
    tmp(36977) := x"0967";
    tmp(36978) := x"0967";
    tmp(36979) := x"0987";
    tmp(36980) := x"09a7";
    tmp(36981) := x"0925";
    tmp(36982) := x"00c4";
    tmp(36983) := x"00a3";
    tmp(36984) := x"00e3";
    tmp(36985) := x"0945";
    tmp(36986) := x"0925";
    tmp(36987) := x"08e4";
    tmp(36988) := x"0062";
    tmp(36989) := x"0020";
    tmp(36990) := x"0000";
    tmp(36991) := x"0040";
    tmp(36992) := x"08a1";
    tmp(36993) := x"08e1";
    tmp(36994) := x"1121";
    tmp(36995) := x"1141";
    tmp(36996) := x"1141";
    tmp(36997) := x"1141";
    tmp(36998) := x"1141";
    tmp(36999) := x"1161";
    tmp(37000) := x"1161";
    tmp(37001) := x"1161";
    tmp(37002) := x"1161";
    tmp(37003) := x"1181";
    tmp(37004) := x"1161";
    tmp(37005) := x"1161";
    tmp(37006) := x"1161";
    tmp(37007) := x"1140";
    tmp(37008) := x"1140";
    tmp(37009) := x"1140";
    tmp(37010) := x"0920";
    tmp(37011) := x"1120";
    tmp(37012) := x"1140";
    tmp(37013) := x"1140";
    tmp(37014) := x"1140";
    tmp(37015) := x"1140";
    tmp(37016) := x"1160";
    tmp(37017) := x"1140";
    tmp(37018) := x"1160";
    tmp(37019) := x"1160";
    tmp(37020) := x"1140";
    tmp(37021) := x"1140";
    tmp(37022) := x"1140";
    tmp(37023) := x"1140";
    tmp(37024) := x"1140";
    tmp(37025) := x"1161";
    tmp(37026) := x"1140";
    tmp(37027) := x"1140";
    tmp(37028) := x"1140";
    tmp(37029) := x"1141";
    tmp(37030) := x"1140";
    tmp(37031) := x"1140";
    tmp(37032) := x"1140";
    tmp(37033) := x"1120";
    tmp(37034) := x"1120";
    tmp(37035) := x"1120";
    tmp(37036) := x"0920";
    tmp(37037) := x"0920";
    tmp(37038) := x"0920";
    tmp(37039) := x"0900";
    tmp(37040) := x"0920";
    tmp(37041) := x"0900";
    tmp(37042) := x"0900";
    tmp(37043) := x"0900";
    tmp(37044) := x"1121";
    tmp(37045) := x"1121";
    tmp(37046) := x"1121";
    tmp(37047) := x"1121";
    tmp(37048) := x"1121";
    tmp(37049) := x"1121";
    tmp(37050) := x"1101";
    tmp(37051) := x"1121";
    tmp(37052) := x"1121";
    tmp(37053) := x"1121";
    tmp(37054) := x"1121";
    tmp(37055) := x"1141";
    tmp(37056) := x"1941";
    tmp(37057) := x"1941";
    tmp(37058) := x"1141";
    tmp(37059) := x"1141";
    tmp(37060) := x"1141";
    tmp(37061) := x"1121";
    tmp(37062) := x"1121";
    tmp(37063) := x"0900";
    tmp(37064) := x"0900";
    tmp(37065) := x"08e0";
    tmp(37066) := x"08e0";
    tmp(37067) := x"0900";
    tmp(37068) := x"08e0";
    tmp(37069) := x"08e0";
    tmp(37070) := x"08e0";
    tmp(37071) := x"08e0";
    tmp(37072) := x"08e0";
    tmp(37073) := x"08e0";
    tmp(37074) := x"08e0";
    tmp(37075) := x"08c0";
    tmp(37076) := x"08e0";
    tmp(37077) := x"10e0";
    tmp(37078) := x"10e0";
    tmp(37079) := x"10e0";
    tmp(37080) := x"1100";
    tmp(37081) := x"10e0";
    tmp(37082) := x"08c0";
    tmp(37083) := x"08c0";
    tmp(37084) := x"08c0";
    tmp(37085) := x"08c0";
    tmp(37086) := x"08e0";
    tmp(37087) := x"08e0";
    tmp(37088) := x"08e0";
    tmp(37089) := x"08e0";
    tmp(37090) := x"0900";
    tmp(37091) := x"0900";
    tmp(37092) := x"0900";
    tmp(37093) := x"0900";
    tmp(37094) := x"0900";
    tmp(37095) := x"0900";
    tmp(37096) := x"0900";
    tmp(37097) := x"0900";
    tmp(37098) := x"08e0";
    tmp(37099) := x"08e0";
    tmp(37100) := x"08e0";
    tmp(37101) := x"08e0";
    tmp(37102) := x"08c0";
    tmp(37103) := x"08c0";
    tmp(37104) := x"08c0";
    tmp(37105) := x"08a0";
    tmp(37106) := x"08a0";
    tmp(37107) := x"08a0";
    tmp(37108) := x"08a0";
    tmp(37109) := x"0880";
    tmp(37110) := x"0880";
    tmp(37111) := x"0880";
    tmp(37112) := x"0880";
    tmp(37113) := x"1080";
    tmp(37114) := x"0880";
    tmp(37115) := x"1080";
    tmp(37116) := x"1080";
    tmp(37117) := x"1080";
    tmp(37118) := x"1060";
    tmp(37119) := x"1060";
    tmp(37120) := x"1060";
    tmp(37121) := x"1060";
    tmp(37122) := x"1060";
    tmp(37123) := x"1060";
    tmp(37124) := x"1060";
    tmp(37125) := x"1060";
    tmp(37126) := x"1060";
    tmp(37127) := x"1060";
    tmp(37128) := x"1060";
    tmp(37129) := x"1040";
    tmp(37130) := x"1040";
    tmp(37131) := x"1040";
    tmp(37132) := x"1040";
    tmp(37133) := x"1040";
    tmp(37134) := x"1040";
    tmp(37135) := x"1040";
    tmp(37136) := x"1060";
    tmp(37137) := x"1060";
    tmp(37138) := x"1060";
    tmp(37139) := x"1060";
    tmp(37140) := x"1060";
    tmp(37141) := x"1060";
    tmp(37142) := x"1061";
    tmp(37143) := x"1061";
    tmp(37144) := x"1060";
    tmp(37145) := x"1060";
    tmp(37146) := x"1060";
    tmp(37147) := x"1060";
    tmp(37148) := x"1060";
    tmp(37149) := x"1060";
    tmp(37150) := x"1060";
    tmp(37151) := x"1040";
    tmp(37152) := x"1040";
    tmp(37153) := x"1040";
    tmp(37154) := x"1040";
    tmp(37155) := x"1040";
    tmp(37156) := x"1040";
    tmp(37157) := x"07e0";
    tmp(37158) := x"07e0";
    tmp(37159) := x"07e0";
    tmp(37160) := x"07e0";
    tmp(37161) := x"07e0";
    tmp(37162) := x"07e0";
    tmp(37163) := x"07e0";
    tmp(37164) := x"07e0";
    tmp(37165) := x"07e0";
    tmp(37166) := x"07e0";
    tmp(37167) := x"07e0";
    tmp(37168) := x"07e0";
    tmp(37169) := x"07e0";
    tmp(37170) := x"07e0";
    tmp(37171) := x"07e0";
    tmp(37172) := x"07e0";
    tmp(37173) := x"07e0";
    tmp(37174) := x"07e0";
    tmp(37175) := x"07e0";
    tmp(37176) := x"07e0";
    tmp(37177) := x"07e0";
    tmp(37178) := x"07e0";
    tmp(37179) := x"07e0";
    tmp(37180) := x"07e0";
    tmp(37181) := x"07e0";
    tmp(37182) := x"07e0";
    tmp(37183) := x"07e0";
    tmp(37184) := x"07e0";
    tmp(37185) := x"07e0";
    tmp(37186) := x"07e0";
    tmp(37187) := x"07e0";
    tmp(37188) := x"07e0";
    tmp(37189) := x"07e0";
    tmp(37190) := x"07e0";
    tmp(37191) := x"07e0";
    tmp(37192) := x"07e0";
    tmp(37193) := x"07e0";
    tmp(37194) := x"07e0";
    tmp(37195) := x"07e0";
    tmp(37196) := x"07e0";
    tmp(37197) := x"0840";
    tmp(37198) := x"0840";
    tmp(37199) := x"0840";
    tmp(37200) := x"0020";
    tmp(37201) := x"0926";
    tmp(37202) := x"0947";
    tmp(37203) := x"0988";
    tmp(37204) := x"0967";
    tmp(37205) := x"0946";
    tmp(37206) := x"0967";
    tmp(37207) := x"0988";
    tmp(37208) := x"0947";
    tmp(37209) := x"0967";
    tmp(37210) := x"09a9";
    tmp(37211) := x"0988";
    tmp(37212) := x"0947";
    tmp(37213) := x"0968";
    tmp(37214) := x"0988";
    tmp(37215) := x"09a8";
    tmp(37216) := x"09e9";
    tmp(37217) := x"122a";
    tmp(37218) := x"11e8";
    tmp(37219) := x"0904";
    tmp(37220) := x"0061";
    tmp(37221) := x"0020";
    tmp(37222) := x"0061";
    tmp(37223) := x"0904";
    tmp(37224) := x"09c7";
    tmp(37225) := x"0904";
    tmp(37226) := x"0041";
    tmp(37227) := x"0000";
    tmp(37228) := x"0000";
    tmp(37229) := x"0020";
    tmp(37230) := x"0880";
    tmp(37231) := x"1101";
    tmp(37232) := x"1141";
    tmp(37233) := x"1121";
    tmp(37234) := x"1120";
    tmp(37235) := x"1120";
    tmp(37236) := x"1120";
    tmp(37237) := x"1141";
    tmp(37238) := x"1161";
    tmp(37239) := x"1161";
    tmp(37240) := x"1161";
    tmp(37241) := x"1161";
    tmp(37242) := x"1181";
    tmp(37243) := x"1181";
    tmp(37244) := x"1181";
    tmp(37245) := x"1181";
    tmp(37246) := x"1161";
    tmp(37247) := x"1160";
    tmp(37248) := x"1140";
    tmp(37249) := x"1140";
    tmp(37250) := x"1140";
    tmp(37251) := x"1140";
    tmp(37252) := x"1140";
    tmp(37253) := x"1140";
    tmp(37254) := x"1160";
    tmp(37255) := x"1140";
    tmp(37256) := x"1160";
    tmp(37257) := x"1140";
    tmp(37258) := x"1140";
    tmp(37259) := x"1140";
    tmp(37260) := x"1141";
    tmp(37261) := x"1140";
    tmp(37262) := x"1140";
    tmp(37263) := x"1140";
    tmp(37264) := x"1140";
    tmp(37265) := x"1161";
    tmp(37266) := x"1160";
    tmp(37267) := x"1141";
    tmp(37268) := x"1141";
    tmp(37269) := x"1141";
    tmp(37270) := x"1140";
    tmp(37271) := x"1140";
    tmp(37272) := x"1140";
    tmp(37273) := x"1120";
    tmp(37274) := x"1120";
    tmp(37275) := x"0920";
    tmp(37276) := x"0920";
    tmp(37277) := x"0920";
    tmp(37278) := x"0920";
    tmp(37279) := x"0920";
    tmp(37280) := x"0920";
    tmp(37281) := x"0900";
    tmp(37282) := x"0900";
    tmp(37283) := x"0900";
    tmp(37284) := x"0900";
    tmp(37285) := x"1120";
    tmp(37286) := x"1121";
    tmp(37287) := x"1121";
    tmp(37288) := x"1121";
    tmp(37289) := x"1121";
    tmp(37290) := x"1101";
    tmp(37291) := x"1121";
    tmp(37292) := x"1121";
    tmp(37293) := x"1121";
    tmp(37294) := x"1141";
    tmp(37295) := x"1141";
    tmp(37296) := x"1141";
    tmp(37297) := x"1141";
    tmp(37298) := x"1141";
    tmp(37299) := x"1141";
    tmp(37300) := x"1121";
    tmp(37301) := x"1121";
    tmp(37302) := x"1121";
    tmp(37303) := x"0900";
    tmp(37304) := x"0900";
    tmp(37305) := x"0900";
    tmp(37306) := x"0900";
    tmp(37307) := x"0900";
    tmp(37308) := x"08e0";
    tmp(37309) := x"08e0";
    tmp(37310) := x"08e0";
    tmp(37311) := x"08e0";
    tmp(37312) := x"08e0";
    tmp(37313) := x"08c0";
    tmp(37314) := x"08e0";
    tmp(37315) := x"08e0";
    tmp(37316) := x"08e0";
    tmp(37317) := x"10e0";
    tmp(37318) := x"10e0";
    tmp(37319) := x"1100";
    tmp(37320) := x"10e0";
    tmp(37321) := x"10e0";
    tmp(37322) := x"08c0";
    tmp(37323) := x"08c0";
    tmp(37324) := x"08c0";
    tmp(37325) := x"08c0";
    tmp(37326) := x"08c0";
    tmp(37327) := x"08e0";
    tmp(37328) := x"08e0";
    tmp(37329) := x"08e0";
    tmp(37330) := x"08e0";
    tmp(37331) := x"0900";
    tmp(37332) := x"0900";
    tmp(37333) := x"0900";
    tmp(37334) := x"0900";
    tmp(37335) := x"0900";
    tmp(37336) := x"0900";
    tmp(37337) := x"0900";
    tmp(37338) := x"0900";
    tmp(37339) := x"08e0";
    tmp(37340) := x"08e0";
    tmp(37341) := x"08c0";
    tmp(37342) := x"08c0";
    tmp(37343) := x"08c0";
    tmp(37344) := x"08c0";
    tmp(37345) := x"08c0";
    tmp(37346) := x"08a0";
    tmp(37347) := x"08a0";
    tmp(37348) := x"0880";
    tmp(37349) := x"1080";
    tmp(37350) := x"1080";
    tmp(37351) := x"1080";
    tmp(37352) := x"1080";
    tmp(37353) := x"1080";
    tmp(37354) := x"1080";
    tmp(37355) := x"1080";
    tmp(37356) := x"1080";
    tmp(37357) := x"1060";
    tmp(37358) := x"1060";
    tmp(37359) := x"1060";
    tmp(37360) := x"1060";
    tmp(37361) := x"1060";
    tmp(37362) := x"1060";
    tmp(37363) := x"1060";
    tmp(37364) := x"1060";
    tmp(37365) := x"1060";
    tmp(37366) := x"1060";
    tmp(37367) := x"1060";
    tmp(37368) := x"1060";
    tmp(37369) := x"1060";
    tmp(37370) := x"1040";
    tmp(37371) := x"1040";
    tmp(37372) := x"1040";
    tmp(37373) := x"1040";
    tmp(37374) := x"1060";
    tmp(37375) := x"1040";
    tmp(37376) := x"1060";
    tmp(37377) := x"1060";
    tmp(37378) := x"1060";
    tmp(37379) := x"1060";
    tmp(37380) := x"1060";
    tmp(37381) := x"1060";
    tmp(37382) := x"1061";
    tmp(37383) := x"1061";
    tmp(37384) := x"1061";
    tmp(37385) := x"1060";
    tmp(37386) := x"1061";
    tmp(37387) := x"1060";
    tmp(37388) := x"1060";
    tmp(37389) := x"1060";
    tmp(37390) := x"1060";
    tmp(37391) := x"1040";
    tmp(37392) := x"1060";
    tmp(37393) := x"1040";
    tmp(37394) := x"1040";
    tmp(37395) := x"1040";
    tmp(37396) := x"1040";
    tmp(37397) := x"07e0";
    tmp(37398) := x"07e0";
    tmp(37399) := x"07e0";
    tmp(37400) := x"07e0";
    tmp(37401) := x"07e0";
    tmp(37402) := x"07e0";
    tmp(37403) := x"07e0";
    tmp(37404) := x"07e0";
    tmp(37405) := x"07e0";
    tmp(37406) := x"07e0";
    tmp(37407) := x"07e0";
    tmp(37408) := x"07e0";
    tmp(37409) := x"07e0";
    tmp(37410) := x"07e0";
    tmp(37411) := x"07e0";
    tmp(37412) := x"07e0";
    tmp(37413) := x"07e0";
    tmp(37414) := x"07e0";
    tmp(37415) := x"07e0";
    tmp(37416) := x"07e0";
    tmp(37417) := x"07e0";
    tmp(37418) := x"07e0";
    tmp(37419) := x"07e0";
    tmp(37420) := x"07e0";
    tmp(37421) := x"07e0";
    tmp(37422) := x"07e0";
    tmp(37423) := x"07e0";
    tmp(37424) := x"07e0";
    tmp(37425) := x"07e0";
    tmp(37426) := x"07e0";
    tmp(37427) := x"07e0";
    tmp(37428) := x"07e0";
    tmp(37429) := x"07e0";
    tmp(37430) := x"07e0";
    tmp(37431) := x"07e0";
    tmp(37432) := x"07e0";
    tmp(37433) := x"07e0";
    tmp(37434) := x"07e0";
    tmp(37435) := x"07e0";
    tmp(37436) := x"07e0";
    tmp(37437) := x"0840";
    tmp(37438) := x"0840";
    tmp(37439) := x"0840";
    tmp(37440) := x"0021";
    tmp(37441) := x"0988";
    tmp(37442) := x"09c9";
    tmp(37443) := x"09a8";
    tmp(37444) := x"0988";
    tmp(37445) := x"0988";
    tmp(37446) := x"09ea";
    tmp(37447) := x"0a0a";
    tmp(37448) := x"09ca";
    tmp(37449) := x"09ca";
    tmp(37450) := x"0967";
    tmp(37451) := x"0947";
    tmp(37452) := x"09a9";
    tmp(37453) := x"0a0a";
    tmp(37454) := x"0a4b";
    tmp(37455) := x"126b";
    tmp(37456) := x"09c7";
    tmp(37457) := x"08c3";
    tmp(37458) := x"0041";
    tmp(37459) := x"0020";
    tmp(37460) := x"0040";
    tmp(37461) := x"0903";
    tmp(37462) := x"1249";
    tmp(37463) := x"09a7";
    tmp(37464) := x"0081";
    tmp(37465) := x"0020";
    tmp(37466) := x"0000";
    tmp(37467) := x"0020";
    tmp(37468) := x"0860";
    tmp(37469) := x"08c1";
    tmp(37470) := x"1121";
    tmp(37471) := x"1141";
    tmp(37472) := x"1141";
    tmp(37473) := x"1120";
    tmp(37474) := x"1121";
    tmp(37475) := x"1120";
    tmp(37476) := x"1140";
    tmp(37477) := x"1141";
    tmp(37478) := x"1161";
    tmp(37479) := x"1161";
    tmp(37480) := x"1181";
    tmp(37481) := x"1181";
    tmp(37482) := x"1181";
    tmp(37483) := x"1181";
    tmp(37484) := x"1161";
    tmp(37485) := x"1181";
    tmp(37486) := x"1181";
    tmp(37487) := x"1161";
    tmp(37488) := x"1160";
    tmp(37489) := x"1140";
    tmp(37490) := x"1140";
    tmp(37491) := x"1140";
    tmp(37492) := x"1140";
    tmp(37493) := x"1140";
    tmp(37494) := x"1140";
    tmp(37495) := x"1160";
    tmp(37496) := x"1161";
    tmp(37497) := x"1160";
    tmp(37498) := x"1161";
    tmp(37499) := x"1140";
    tmp(37500) := x"1160";
    tmp(37501) := x"1160";
    tmp(37502) := x"1140";
    tmp(37503) := x"1141";
    tmp(37504) := x"1160";
    tmp(37505) := x"1141";
    tmp(37506) := x"1141";
    tmp(37507) := x"1141";
    tmp(37508) := x"1141";
    tmp(37509) := x"1141";
    tmp(37510) := x"1141";
    tmp(37511) := x"1120";
    tmp(37512) := x"1141";
    tmp(37513) := x"1140";
    tmp(37514) := x"1140";
    tmp(37515) := x"1120";
    tmp(37516) := x"1120";
    tmp(37517) := x"1120";
    tmp(37518) := x"0920";
    tmp(37519) := x"0920";
    tmp(37520) := x"0920";
    tmp(37521) := x"0920";
    tmp(37522) := x"0900";
    tmp(37523) := x"0900";
    tmp(37524) := x"0900";
    tmp(37525) := x"0900";
    tmp(37526) := x"1120";
    tmp(37527) := x"1121";
    tmp(37528) := x"1121";
    tmp(37529) := x"1121";
    tmp(37530) := x"1121";
    tmp(37531) := x"1121";
    tmp(37532) := x"1141";
    tmp(37533) := x"1141";
    tmp(37534) := x"1141";
    tmp(37535) := x"1141";
    tmp(37536) := x"1141";
    tmp(37537) := x"1141";
    tmp(37538) := x"1141";
    tmp(37539) := x"1141";
    tmp(37540) := x"1121";
    tmp(37541) := x"1121";
    tmp(37542) := x"0900";
    tmp(37543) := x"0900";
    tmp(37544) := x"0900";
    tmp(37545) := x"0900";
    tmp(37546) := x"0900";
    tmp(37547) := x"08e0";
    tmp(37548) := x"0900";
    tmp(37549) := x"08e0";
    tmp(37550) := x"08e0";
    tmp(37551) := x"08e0";
    tmp(37552) := x"08c0";
    tmp(37553) := x"08e0";
    tmp(37554) := x"08c0";
    tmp(37555) := x"08e0";
    tmp(37556) := x"08e0";
    tmp(37557) := x"08e0";
    tmp(37558) := x"10e0";
    tmp(37559) := x"1100";
    tmp(37560) := x"10e0";
    tmp(37561) := x"10e0";
    tmp(37562) := x"08c0";
    tmp(37563) := x"08c0";
    tmp(37564) := x"08c0";
    tmp(37565) := x"08c0";
    tmp(37566) := x"08c0";
    tmp(37567) := x"08e0";
    tmp(37568) := x"08e0";
    tmp(37569) := x"08e0";
    tmp(37570) := x"08e0";
    tmp(37571) := x"0900";
    tmp(37572) := x"0900";
    tmp(37573) := x"0900";
    tmp(37574) := x"0900";
    tmp(37575) := x"0900";
    tmp(37576) := x"0900";
    tmp(37577) := x"0900";
    tmp(37578) := x"0900";
    tmp(37579) := x"0900";
    tmp(37580) := x"08e0";
    tmp(37581) := x"08e0";
    tmp(37582) := x"08c0";
    tmp(37583) := x"08c0";
    tmp(37584) := x"08c0";
    tmp(37585) := x"08c0";
    tmp(37586) := x"08a0";
    tmp(37587) := x"08a0";
    tmp(37588) := x"08a0";
    tmp(37589) := x"1080";
    tmp(37590) := x"1080";
    tmp(37591) := x"1080";
    tmp(37592) := x"1080";
    tmp(37593) := x"1080";
    tmp(37594) := x"1080";
    tmp(37595) := x"1080";
    tmp(37596) := x"1080";
    tmp(37597) := x"1060";
    tmp(37598) := x"1060";
    tmp(37599) := x"1060";
    tmp(37600) := x"1060";
    tmp(37601) := x"1060";
    tmp(37602) := x"1060";
    tmp(37603) := x"1060";
    tmp(37604) := x"1060";
    tmp(37605) := x"1060";
    tmp(37606) := x"1060";
    tmp(37607) := x"1060";
    tmp(37608) := x"1060";
    tmp(37609) := x"1060";
    tmp(37610) := x"1040";
    tmp(37611) := x"1040";
    tmp(37612) := x"1040";
    tmp(37613) := x"1040";
    tmp(37614) := x"1060";
    tmp(37615) := x"1040";
    tmp(37616) := x"1040";
    tmp(37617) := x"1060";
    tmp(37618) := x"1060";
    tmp(37619) := x"1060";
    tmp(37620) := x"1060";
    tmp(37621) := x"1060";
    tmp(37622) := x"1061";
    tmp(37623) := x"1061";
    tmp(37624) := x"1061";
    tmp(37625) := x"1061";
    tmp(37626) := x"1061";
    tmp(37627) := x"1061";
    tmp(37628) := x"1061";
    tmp(37629) := x"1061";
    tmp(37630) := x"1060";
    tmp(37631) := x"1060";
    tmp(37632) := x"1040";
    tmp(37633) := x"1040";
    tmp(37634) := x"1040";
    tmp(37635) := x"1060";
    tmp(37636) := x"1040";
    tmp(37637) := x"07e0";
    tmp(37638) := x"07e0";
    tmp(37639) := x"07e0";
    tmp(37640) := x"07e0";
    tmp(37641) := x"07e0";
    tmp(37642) := x"07e0";
    tmp(37643) := x"07e0";
    tmp(37644) := x"07e0";
    tmp(37645) := x"07e0";
    tmp(37646) := x"07e0";
    tmp(37647) := x"07e0";
    tmp(37648) := x"07e0";
    tmp(37649) := x"07e0";
    tmp(37650) := x"07e0";
    tmp(37651) := x"07e0";
    tmp(37652) := x"07e0";
    tmp(37653) := x"07e0";
    tmp(37654) := x"07e0";
    tmp(37655) := x"07e0";
    tmp(37656) := x"07e0";
    tmp(37657) := x"07e0";
    tmp(37658) := x"07e0";
    tmp(37659) := x"07e0";
    tmp(37660) := x"07e0";
    tmp(37661) := x"07e0";
    tmp(37662) := x"07e0";
    tmp(37663) := x"07e0";
    tmp(37664) := x"07e0";
    tmp(37665) := x"07e0";
    tmp(37666) := x"07e0";
    tmp(37667) := x"07e0";
    tmp(37668) := x"07e0";
    tmp(37669) := x"07e0";
    tmp(37670) := x"07e0";
    tmp(37671) := x"07e0";
    tmp(37672) := x"07e0";
    tmp(37673) := x"07e0";
    tmp(37674) := x"07e0";
    tmp(37675) := x"07e0";
    tmp(37676) := x"07e0";
    tmp(37677) := x"1060";
    tmp(37678) := x"0840";
    tmp(37679) := x"0860";
    tmp(37680) := x"0021";
    tmp(37681) := x"09a9";
    tmp(37682) := x"0988";
    tmp(37683) := x"0926";
    tmp(37684) := x"0988";
    tmp(37685) := x"09ea";
    tmp(37686) := x"0a2b";
    tmp(37687) := x"0a2b";
    tmp(37688) := x"0a2b";
    tmp(37689) := x"0988";
    tmp(37690) := x"0926";
    tmp(37691) := x"0987";
    tmp(37692) := x"09a9";
    tmp(37693) := x"09a7";
    tmp(37694) := x"00c3";
    tmp(37695) := x"0041";
    tmp(37696) := x"0020";
    tmp(37697) := x"0000";
    tmp(37698) := x"0020";
    tmp(37699) := x"08c2";
    tmp(37700) := x"1249";
    tmp(37701) := x"126a";
    tmp(37702) := x"0903";
    tmp(37703) := x"0061";
    tmp(37704) := x"0040";
    tmp(37705) := x"0860";
    tmp(37706) := x"08c1";
    tmp(37707) := x"08e1";
    tmp(37708) := x"1101";
    tmp(37709) := x"1120";
    tmp(37710) := x"1120";
    tmp(37711) := x"1140";
    tmp(37712) := x"1141";
    tmp(37713) := x"1141";
    tmp(37714) := x"1121";
    tmp(37715) := x"1120";
    tmp(37716) := x"1141";
    tmp(37717) := x"1141";
    tmp(37718) := x"1161";
    tmp(37719) := x"1181";
    tmp(37720) := x"1181";
    tmp(37721) := x"1161";
    tmp(37722) := x"1181";
    tmp(37723) := x"1161";
    tmp(37724) := x"1161";
    tmp(37725) := x"1981";
    tmp(37726) := x"19a1";
    tmp(37727) := x"1161";
    tmp(37728) := x"1161";
    tmp(37729) := x"1160";
    tmp(37730) := x"1160";
    tmp(37731) := x"1160";
    tmp(37732) := x"1160";
    tmp(37733) := x"1161";
    tmp(37734) := x"1140";
    tmp(37735) := x"1161";
    tmp(37736) := x"1161";
    tmp(37737) := x"1160";
    tmp(37738) := x"1161";
    tmp(37739) := x"1140";
    tmp(37740) := x"1161";
    tmp(37741) := x"1161";
    tmp(37742) := x"1161";
    tmp(37743) := x"1140";
    tmp(37744) := x"1140";
    tmp(37745) := x"1140";
    tmp(37746) := x"1141";
    tmp(37747) := x"1141";
    tmp(37748) := x"1140";
    tmp(37749) := x"1140";
    tmp(37750) := x"1141";
    tmp(37751) := x"1140";
    tmp(37752) := x"1141";
    tmp(37753) := x"1141";
    tmp(37754) := x"1140";
    tmp(37755) := x"1140";
    tmp(37756) := x"1120";
    tmp(37757) := x"0920";
    tmp(37758) := x"0920";
    tmp(37759) := x"0920";
    tmp(37760) := x"0920";
    tmp(37761) := x"0920";
    tmp(37762) := x"0920";
    tmp(37763) := x"0900";
    tmp(37764) := x"0900";
    tmp(37765) := x"0900";
    tmp(37766) := x"0920";
    tmp(37767) := x"0920";
    tmp(37768) := x"0900";
    tmp(37769) := x"1121";
    tmp(37770) := x"1121";
    tmp(37771) := x"1121";
    tmp(37772) := x"1121";
    tmp(37773) := x"1141";
    tmp(37774) := x"1141";
    tmp(37775) := x"1141";
    tmp(37776) := x"1141";
    tmp(37777) := x"1141";
    tmp(37778) := x"1141";
    tmp(37779) := x"1121";
    tmp(37780) := x"1121";
    tmp(37781) := x"0921";
    tmp(37782) := x"0900";
    tmp(37783) := x"0900";
    tmp(37784) := x"0900";
    tmp(37785) := x"0900";
    tmp(37786) := x"0900";
    tmp(37787) := x"0900";
    tmp(37788) := x"0900";
    tmp(37789) := x"08e0";
    tmp(37790) := x"08e0";
    tmp(37791) := x"08e0";
    tmp(37792) := x"08c0";
    tmp(37793) := x"08e0";
    tmp(37794) := x"08e0";
    tmp(37795) := x"08e0";
    tmp(37796) := x"08e0";
    tmp(37797) := x"10e0";
    tmp(37798) := x"10e0";
    tmp(37799) := x"10e0";
    tmp(37800) := x"08e0";
    tmp(37801) := x"08e0";
    tmp(37802) := x"08c0";
    tmp(37803) := x"08c0";
    tmp(37804) := x"08c0";
    tmp(37805) := x"08c0";
    tmp(37806) := x"08c0";
    tmp(37807) := x"08c0";
    tmp(37808) := x"08e0";
    tmp(37809) := x"08e0";
    tmp(37810) := x"08e0";
    tmp(37811) := x"08e0";
    tmp(37812) := x"0900";
    tmp(37813) := x"0900";
    tmp(37814) := x"0900";
    tmp(37815) := x"0900";
    tmp(37816) := x"0900";
    tmp(37817) := x"0900";
    tmp(37818) := x"0900";
    tmp(37819) := x"08e0";
    tmp(37820) := x"08e0";
    tmp(37821) := x"08e0";
    tmp(37822) := x"08e0";
    tmp(37823) := x"08c0";
    tmp(37824) := x"08c0";
    tmp(37825) := x"08c0";
    tmp(37826) := x"08a0";
    tmp(37827) := x"10a0";
    tmp(37828) := x"08a0";
    tmp(37829) := x"1080";
    tmp(37830) := x"1080";
    tmp(37831) := x"1080";
    tmp(37832) := x"1080";
    tmp(37833) := x"1080";
    tmp(37834) := x"1080";
    tmp(37835) := x"1080";
    tmp(37836) := x"1080";
    tmp(37837) := x"1060";
    tmp(37838) := x"1060";
    tmp(37839) := x"1060";
    tmp(37840) := x"1060";
    tmp(37841) := x"1060";
    tmp(37842) := x"1060";
    tmp(37843) := x"1060";
    tmp(37844) := x"1060";
    tmp(37845) := x"1060";
    tmp(37846) := x"1060";
    tmp(37847) := x"1060";
    tmp(37848) := x"1060";
    tmp(37849) := x"1040";
    tmp(37850) := x"1040";
    tmp(37851) := x"1040";
    tmp(37852) := x"1040";
    tmp(37853) := x"1040";
    tmp(37854) := x"1040";
    tmp(37855) := x"1040";
    tmp(37856) := x"1060";
    tmp(37857) := x"1060";
    tmp(37858) := x"1060";
    tmp(37859) := x"1061";
    tmp(37860) := x"1061";
    tmp(37861) := x"1061";
    tmp(37862) := x"1061";
    tmp(37863) := x"1061";
    tmp(37864) := x"1061";
    tmp(37865) := x"1061";
    tmp(37866) := x"1061";
    tmp(37867) := x"1060";
    tmp(37868) := x"1061";
    tmp(37869) := x"1061";
    tmp(37870) := x"1060";
    tmp(37871) := x"1060";
    tmp(37872) := x"1040";
    tmp(37873) := x"1060";
    tmp(37874) := x"1060";
    tmp(37875) := x"1040";
    tmp(37876) := x"1060";
    tmp(37877) := x"07e0";
    tmp(37878) := x"07e0";
    tmp(37879) := x"07e0";
    tmp(37880) := x"07e0";
    tmp(37881) := x"07e0";
    tmp(37882) := x"07e0";
    tmp(37883) := x"07e0";
    tmp(37884) := x"07e0";
    tmp(37885) := x"07e0";
    tmp(37886) := x"07e0";
    tmp(37887) := x"07e0";
    tmp(37888) := x"07e0";
    tmp(37889) := x"07e0";
    tmp(37890) := x"07e0";
    tmp(37891) := x"07e0";
    tmp(37892) := x"07e0";
    tmp(37893) := x"07e0";
    tmp(37894) := x"07e0";
    tmp(37895) := x"07e0";
    tmp(37896) := x"07e0";
    tmp(37897) := x"07e0";
    tmp(37898) := x"07e0";
    tmp(37899) := x"07e0";
    tmp(37900) := x"07e0";
    tmp(37901) := x"07e0";
    tmp(37902) := x"07e0";
    tmp(37903) := x"07e0";
    tmp(37904) := x"07e0";
    tmp(37905) := x"07e0";
    tmp(37906) := x"07e0";
    tmp(37907) := x"07e0";
    tmp(37908) := x"07e0";
    tmp(37909) := x"07e0";
    tmp(37910) := x"07e0";
    tmp(37911) := x"07e0";
    tmp(37912) := x"07e0";
    tmp(37913) := x"07e0";
    tmp(37914) := x"07e0";
    tmp(37915) := x"07e0";
    tmp(37916) := x"07e0";
    tmp(37917) := x"0840";
    tmp(37918) := x"1060";
    tmp(37919) := x"1060";
    tmp(37920) := x"0021";
    tmp(37921) := x"09a9";
    tmp(37922) := x"0967";
    tmp(37923) := x"0967";
    tmp(37924) := x"09ea";
    tmp(37925) := x"0a0a";
    tmp(37926) := x"09ea";
    tmp(37927) := x"09a9";
    tmp(37928) := x"0988";
    tmp(37929) := x"08e5";
    tmp(37930) := x"00c4";
    tmp(37931) := x"00a2";
    tmp(37932) := x"0041";
    tmp(37933) := x"0020";
    tmp(37934) := x"0000";
    tmp(37935) := x"0000";
    tmp(37936) := x"0020";
    tmp(37937) := x"08c2";
    tmp(37938) := x"0986";
    tmp(37939) := x"11e8";
    tmp(37940) := x"0924";
    tmp(37941) := x"08c1";
    tmp(37942) := x"08e1";
    tmp(37943) := x"0901";
    tmp(37944) := x"1121";
    tmp(37945) := x"1121";
    tmp(37946) := x"1141";
    tmp(37947) := x"1121";
    tmp(37948) := x"1120";
    tmp(37949) := x"1120";
    tmp(37950) := x"1120";
    tmp(37951) := x"1140";
    tmp(37952) := x"1141";
    tmp(37953) := x"1141";
    tmp(37954) := x"1141";
    tmp(37955) := x"1141";
    tmp(37956) := x"1141";
    tmp(37957) := x"1141";
    tmp(37958) := x"1161";
    tmp(37959) := x"1181";
    tmp(37960) := x"1181";
    tmp(37961) := x"1981";
    tmp(37962) := x"1981";
    tmp(37963) := x"1181";
    tmp(37964) := x"1161";
    tmp(37965) := x"1981";
    tmp(37966) := x"1981";
    tmp(37967) := x"1181";
    tmp(37968) := x"1181";
    tmp(37969) := x"1161";
    tmp(37970) := x"1161";
    tmp(37971) := x"1161";
    tmp(37972) := x"1160";
    tmp(37973) := x"1161";
    tmp(37974) := x"1161";
    tmp(37975) := x"1161";
    tmp(37976) := x"1181";
    tmp(37977) := x"1161";
    tmp(37978) := x"1161";
    tmp(37979) := x"1141";
    tmp(37980) := x"1141";
    tmp(37981) := x"1161";
    tmp(37982) := x"1141";
    tmp(37983) := x"1140";
    tmp(37984) := x"1161";
    tmp(37985) := x"1141";
    tmp(37986) := x"1141";
    tmp(37987) := x"1141";
    tmp(37988) := x"1140";
    tmp(37989) := x"1140";
    tmp(37990) := x"1140";
    tmp(37991) := x"1140";
    tmp(37992) := x"1141";
    tmp(37993) := x"1141";
    tmp(37994) := x"1140";
    tmp(37995) := x"1140";
    tmp(37996) := x"1140";
    tmp(37997) := x"1140";
    tmp(37998) := x"0920";
    tmp(37999) := x"0920";
    tmp(38000) := x"0920";
    tmp(38001) := x"0920";
    tmp(38002) := x"0920";
    tmp(38003) := x"0920";
    tmp(38004) := x"0900";
    tmp(38005) := x"0900";
    tmp(38006) := x"08e0";
    tmp(38007) := x"0900";
    tmp(38008) := x"0920";
    tmp(38009) := x"0920";
    tmp(38010) := x"0920";
    tmp(38011) := x"1121";
    tmp(38012) := x"1141";
    tmp(38013) := x"1121";
    tmp(38014) := x"1121";
    tmp(38015) := x"1141";
    tmp(38016) := x"1141";
    tmp(38017) := x"1141";
    tmp(38018) := x"1141";
    tmp(38019) := x"1121";
    tmp(38020) := x"0921";
    tmp(38021) := x"0900";
    tmp(38022) := x"0900";
    tmp(38023) := x"0900";
    tmp(38024) := x"0900";
    tmp(38025) := x"08e0";
    tmp(38026) := x"08e0";
    tmp(38027) := x"0900";
    tmp(38028) := x"08e0";
    tmp(38029) := x"08e0";
    tmp(38030) := x"08e0";
    tmp(38031) := x"08e0";
    tmp(38032) := x"08e0";
    tmp(38033) := x"08e0";
    tmp(38034) := x"08e0";
    tmp(38035) := x"08e0";
    tmp(38036) := x"08c0";
    tmp(38037) := x"10e0";
    tmp(38038) := x"08e0";
    tmp(38039) := x"08e0";
    tmp(38040) := x"08e0";
    tmp(38041) := x"08e0";
    tmp(38042) := x"08c0";
    tmp(38043) := x"08c0";
    tmp(38044) := x"08c0";
    tmp(38045) := x"08c0";
    tmp(38046) := x"08c0";
    tmp(38047) := x"08c0";
    tmp(38048) := x"08c0";
    tmp(38049) := x"08c0";
    tmp(38050) := x"08c0";
    tmp(38051) := x"08e0";
    tmp(38052) := x"08e0";
    tmp(38053) := x"0900";
    tmp(38054) := x"0900";
    tmp(38055) := x"0900";
    tmp(38056) := x"0900";
    tmp(38057) := x"0900";
    tmp(38058) := x"0900";
    tmp(38059) := x"08e0";
    tmp(38060) := x"08e0";
    tmp(38061) := x"08c0";
    tmp(38062) := x"08c0";
    tmp(38063) := x"08c0";
    tmp(38064) := x"08c0";
    tmp(38065) := x"08c0";
    tmp(38066) := x"08a0";
    tmp(38067) := x"08a0";
    tmp(38068) := x"08a0";
    tmp(38069) := x"1080";
    tmp(38070) := x"1080";
    tmp(38071) := x"0880";
    tmp(38072) := x"1080";
    tmp(38073) := x"1060";
    tmp(38074) := x"1080";
    tmp(38075) := x"1060";
    tmp(38076) := x"1060";
    tmp(38077) := x"1060";
    tmp(38078) := x"1060";
    tmp(38079) := x"1060";
    tmp(38080) := x"1060";
    tmp(38081) := x"1060";
    tmp(38082) := x"1060";
    tmp(38083) := x"1060";
    tmp(38084) := x"1060";
    tmp(38085) := x"1060";
    tmp(38086) := x"1060";
    tmp(38087) := x"1060";
    tmp(38088) := x"1060";
    tmp(38089) := x"1040";
    tmp(38090) := x"1040";
    tmp(38091) := x"1040";
    tmp(38092) := x"1040";
    tmp(38093) := x"1040";
    tmp(38094) := x"1040";
    tmp(38095) := x"1040";
    tmp(38096) := x"1060";
    tmp(38097) := x"1060";
    tmp(38098) := x"1060";
    tmp(38099) := x"1061";
    tmp(38100) := x"1060";
    tmp(38101) := x"1060";
    tmp(38102) := x"1061";
    tmp(38103) := x"1061";
    tmp(38104) := x"1061";
    tmp(38105) := x"1061";
    tmp(38106) := x"1060";
    tmp(38107) := x"1061";
    tmp(38108) := x"1061";
    tmp(38109) := x"1060";
    tmp(38110) := x"1060";
    tmp(38111) := x"1060";
    tmp(38112) := x"1060";
    tmp(38113) := x"1040";
    tmp(38114) := x"1060";
    tmp(38115) := x"1040";
    tmp(38116) := x"1040";
    tmp(38117) := x"07e0";
    tmp(38118) := x"07e0";
    tmp(38119) := x"07e0";
    tmp(38120) := x"07e0";
    tmp(38121) := x"07e0";
    tmp(38122) := x"07e0";
    tmp(38123) := x"07e0";
    tmp(38124) := x"07e0";
    tmp(38125) := x"07e0";
    tmp(38126) := x"07e0";
    tmp(38127) := x"07e0";
    tmp(38128) := x"07e0";
    tmp(38129) := x"07e0";
    tmp(38130) := x"07e0";
    tmp(38131) := x"07e0";
    tmp(38132) := x"07e0";
    tmp(38133) := x"07e0";
    tmp(38134) := x"07e0";
    tmp(38135) := x"07e0";
    tmp(38136) := x"07e0";
    tmp(38137) := x"07e0";
    tmp(38138) := x"07e0";
    tmp(38139) := x"07e0";
    tmp(38140) := x"07e0";
    tmp(38141) := x"07e0";
    tmp(38142) := x"07e0";
    tmp(38143) := x"07e0";
    tmp(38144) := x"07e0";
    tmp(38145) := x"07e0";
    tmp(38146) := x"07e0";
    tmp(38147) := x"07e0";
    tmp(38148) := x"07e0";
    tmp(38149) := x"07e0";
    tmp(38150) := x"07e0";
    tmp(38151) := x"07e0";
    tmp(38152) := x"07e0";
    tmp(38153) := x"07e0";
    tmp(38154) := x"07e0";
    tmp(38155) := x"07e0";
    tmp(38156) := x"07e0";
    tmp(38157) := x"1060";
    tmp(38158) := x"1060";
    tmp(38159) := x"0860";
    tmp(38160) := x"0021";
    tmp(38161) := x"09ca";
    tmp(38162) := x"09a9";
    tmp(38163) := x"09a8";
    tmp(38164) := x"0988";
    tmp(38165) := x"0967";
    tmp(38166) := x"0967";
    tmp(38167) := x"0105";
    tmp(38168) := x"0082";
    tmp(38169) := x"0041";
    tmp(38170) := x"0020";
    tmp(38171) := x"0000";
    tmp(38172) := x"0000";
    tmp(38173) := x"0020";
    tmp(38174) := x"0020";
    tmp(38175) := x"0861";
    tmp(38176) := x"0882";
    tmp(38177) := x"0041";
    tmp(38178) := x"0041";
    tmp(38179) := x"0040";
    tmp(38180) := x"0880";
    tmp(38181) := x"1121";
    tmp(38182) := x"1161";
    tmp(38183) := x"1141";
    tmp(38184) := x"1120";
    tmp(38185) := x"1140";
    tmp(38186) := x"1120";
    tmp(38187) := x"1140";
    tmp(38188) := x"1120";
    tmp(38189) := x"1120";
    tmp(38190) := x"1120";
    tmp(38191) := x"1140";
    tmp(38192) := x"1161";
    tmp(38193) := x"1141";
    tmp(38194) := x"1141";
    tmp(38195) := x"1141";
    tmp(38196) := x"1141";
    tmp(38197) := x"1141";
    tmp(38198) := x"1161";
    tmp(38199) := x"1161";
    tmp(38200) := x"1161";
    tmp(38201) := x"1981";
    tmp(38202) := x"19a1";
    tmp(38203) := x"1981";
    tmp(38204) := x"1181";
    tmp(38205) := x"1981";
    tmp(38206) := x"1181";
    tmp(38207) := x"1181";
    tmp(38208) := x"1181";
    tmp(38209) := x"1181";
    tmp(38210) := x"1161";
    tmp(38211) := x"1161";
    tmp(38212) := x"1161";
    tmp(38213) := x"1161";
    tmp(38214) := x"1161";
    tmp(38215) := x"1181";
    tmp(38216) := x"1181";
    tmp(38217) := x"1181";
    tmp(38218) := x"1160";
    tmp(38219) := x"1160";
    tmp(38220) := x"1161";
    tmp(38221) := x"1161";
    tmp(38222) := x"1140";
    tmp(38223) := x"1141";
    tmp(38224) := x"1140";
    tmp(38225) := x"1140";
    tmp(38226) := x"1140";
    tmp(38227) := x"1141";
    tmp(38228) := x"1161";
    tmp(38229) := x"1161";
    tmp(38230) := x"1140";
    tmp(38231) := x"1140";
    tmp(38232) := x"1141";
    tmp(38233) := x"1161";
    tmp(38234) := x"1140";
    tmp(38235) := x"1141";
    tmp(38236) := x"1120";
    tmp(38237) := x"1141";
    tmp(38238) := x"1140";
    tmp(38239) := x"0940";
    tmp(38240) := x"0920";
    tmp(38241) := x"0920";
    tmp(38242) := x"0920";
    tmp(38243) := x"0900";
    tmp(38244) := x"0900";
    tmp(38245) := x"0900";
    tmp(38246) := x"0900";
    tmp(38247) := x"08e0";
    tmp(38248) := x"0900";
    tmp(38249) := x"0900";
    tmp(38250) := x"0920";
    tmp(38251) := x"0900";
    tmp(38252) := x"1120";
    tmp(38253) := x"1121";
    tmp(38254) := x"1121";
    tmp(38255) := x"1141";
    tmp(38256) := x"1141";
    tmp(38257) := x"1141";
    tmp(38258) := x"1141";
    tmp(38259) := x"0921";
    tmp(38260) := x"0920";
    tmp(38261) := x"0900";
    tmp(38262) := x"0900";
    tmp(38263) := x"0900";
    tmp(38264) := x"08e0";
    tmp(38265) := x"0900";
    tmp(38266) := x"08e0";
    tmp(38267) := x"08e0";
    tmp(38268) := x"08e0";
    tmp(38269) := x"08e0";
    tmp(38270) := x"08e0";
    tmp(38271) := x"08e0";
    tmp(38272) := x"08e0";
    tmp(38273) := x"08e0";
    tmp(38274) := x"08e0";
    tmp(38275) := x"08e0";
    tmp(38276) := x"08e0";
    tmp(38277) := x"08e0";
    tmp(38278) := x"08c0";
    tmp(38279) := x"08c0";
    tmp(38280) := x"08c0";
    tmp(38281) := x"08e0";
    tmp(38282) := x"08e0";
    tmp(38283) := x"08c0";
    tmp(38284) := x"08c0";
    tmp(38285) := x"08c0";
    tmp(38286) := x"08c0";
    tmp(38287) := x"08c0";
    tmp(38288) := x"08c0";
    tmp(38289) := x"08c0";
    tmp(38290) := x"08c0";
    tmp(38291) := x"08c0";
    tmp(38292) := x"08e0";
    tmp(38293) := x"0900";
    tmp(38294) := x"0900";
    tmp(38295) := x"0900";
    tmp(38296) := x"0900";
    tmp(38297) := x"0900";
    tmp(38298) := x"0900";
    tmp(38299) := x"0900";
    tmp(38300) := x"08e0";
    tmp(38301) := x"08e0";
    tmp(38302) := x"08c0";
    tmp(38303) := x"08c0";
    tmp(38304) := x"08c0";
    tmp(38305) := x"08c0";
    tmp(38306) := x"08a0";
    tmp(38307) := x"08a0";
    tmp(38308) := x"0880";
    tmp(38309) := x"1080";
    tmp(38310) := x"1080";
    tmp(38311) := x"1080";
    tmp(38312) := x"1080";
    tmp(38313) := x"1080";
    tmp(38314) := x"1060";
    tmp(38315) := x"1060";
    tmp(38316) := x"1060";
    tmp(38317) := x"1060";
    tmp(38318) := x"1060";
    tmp(38319) := x"1060";
    tmp(38320) := x"1060";
    tmp(38321) := x"1060";
    tmp(38322) := x"1060";
    tmp(38323) := x"1060";
    tmp(38324) := x"1060";
    tmp(38325) := x"1060";
    tmp(38326) := x"1060";
    tmp(38327) := x"1060";
    tmp(38328) := x"1060";
    tmp(38329) := x"1040";
    tmp(38330) := x"1040";
    tmp(38331) := x"1040";
    tmp(38332) := x"1040";
    tmp(38333) := x"1040";
    tmp(38334) := x"1040";
    tmp(38335) := x"1060";
    tmp(38336) := x"1060";
    tmp(38337) := x"1060";
    tmp(38338) := x"1060";
    tmp(38339) := x"1061";
    tmp(38340) := x"1061";
    tmp(38341) := x"1061";
    tmp(38342) := x"1061";
    tmp(38343) := x"1061";
    tmp(38344) := x"1061";
    tmp(38345) := x"1061";
    tmp(38346) := x"1061";
    tmp(38347) := x"1061";
    tmp(38348) := x"1060";
    tmp(38349) := x"1060";
    tmp(38350) := x"1060";
    tmp(38351) := x"1060";
    tmp(38352) := x"1040";
    tmp(38353) := x"1060";
    tmp(38354) := x"1040";
    tmp(38355) := x"1040";
    tmp(38356) := x"1040";
    tmp(38357) := x"07e0";
    tmp(38358) := x"07e0";
    tmp(38359) := x"07e0";
    tmp(38360) := x"07e0";
    tmp(38361) := x"07e0";
    tmp(38362) := x"07e0";
    tmp(38363) := x"07e0";
    tmp(38364) := x"07e0";
    tmp(38365) := x"07e0";
    tmp(38366) := x"07e0";
    tmp(38367) := x"07e0";
    tmp(38368) := x"07e0";
    tmp(38369) := x"07e0";
    tmp(38370) := x"07e0";
    tmp(38371) := x"07e0";
    tmp(38372) := x"07e0";
    tmp(38373) := x"07e0";
    tmp(38374) := x"07e0";
    tmp(38375) := x"07e0";
    tmp(38376) := x"07e0";
    tmp(38377) := x"07e0";
    tmp(38378) := x"07e0";
    tmp(38379) := x"07e0";
    tmp(38380) := x"07e0";
    tmp(38381) := x"07e0";
    tmp(38382) := x"07e0";
    tmp(38383) := x"07e0";
    tmp(38384) := x"07e0";
    tmp(38385) := x"07e0";
    tmp(38386) := x"07e0";
    tmp(38387) := x"07e0";
    tmp(38388) := x"07e0";
    tmp(38389) := x"07e0";
    tmp(38390) := x"07e0";
    tmp(38391) := x"07e0";
    tmp(38392) := x"07e0";
    tmp(38393) := x"07e0";
    tmp(38394) := x"07e0";
    tmp(38395) := x"07e0";
    tmp(38396) := x"07e0";
    tmp(38397) := x"1060";
    tmp(38398) := x"1061";
    tmp(38399) := x"1061";
    tmp(38400) := x"0021";
    tmp(38401) := x"09a8";
    tmp(38402) := x"0967";
    tmp(38403) := x"09a7";
    tmp(38404) := x"09a8";
    tmp(38405) := x"0925";
    tmp(38406) := x"00a3";
    tmp(38407) := x"0062";
    tmp(38408) := x"0021";
    tmp(38409) := x"0041";
    tmp(38410) := x"08c3";
    tmp(38411) := x"08c3";
    tmp(38412) := x"08a2";
    tmp(38413) := x"0061";
    tmp(38414) := x"0020";
    tmp(38415) := x"0000";
    tmp(38416) := x"0000";
    tmp(38417) := x"0020";
    tmp(38418) := x"0040";
    tmp(38419) := x"08c0";
    tmp(38420) := x"1141";
    tmp(38421) := x"1161";
    tmp(38422) := x"1161";
    tmp(38423) := x"1141";
    tmp(38424) := x"1120";
    tmp(38425) := x"1120";
    tmp(38426) := x"1120";
    tmp(38427) := x"1140";
    tmp(38428) := x"1120";
    tmp(38429) := x"1120";
    tmp(38430) := x"1120";
    tmp(38431) := x"1120";
    tmp(38432) := x"1140";
    tmp(38433) := x"1140";
    tmp(38434) := x"1140";
    tmp(38435) := x"1141";
    tmp(38436) := x"1141";
    tmp(38437) := x"1141";
    tmp(38438) := x"1161";
    tmp(38439) := x"1161";
    tmp(38440) := x"1161";
    tmp(38441) := x"1161";
    tmp(38442) := x"1981";
    tmp(38443) := x"1981";
    tmp(38444) := x"19a1";
    tmp(38445) := x"1981";
    tmp(38446) := x"1181";
    tmp(38447) := x"1181";
    tmp(38448) := x"1181";
    tmp(38449) := x"1181";
    tmp(38450) := x"1181";
    tmp(38451) := x"1161";
    tmp(38452) := x"1161";
    tmp(38453) := x"1161";
    tmp(38454) := x"1161";
    tmp(38455) := x"1161";
    tmp(38456) := x"1161";
    tmp(38457) := x"1161";
    tmp(38458) := x"1161";
    tmp(38459) := x"1161";
    tmp(38460) := x"1140";
    tmp(38461) := x"1161";
    tmp(38462) := x"1140";
    tmp(38463) := x"1161";
    tmp(38464) := x"1140";
    tmp(38465) := x"1140";
    tmp(38466) := x"1140";
    tmp(38467) := x"1141";
    tmp(38468) := x"1141";
    tmp(38469) := x"1140";
    tmp(38470) := x"1161";
    tmp(38471) := x"1141";
    tmp(38472) := x"1141";
    tmp(38473) := x"1141";
    tmp(38474) := x"1140";
    tmp(38475) := x"1140";
    tmp(38476) := x"1161";
    tmp(38477) := x"1140";
    tmp(38478) := x"1141";
    tmp(38479) := x"0920";
    tmp(38480) := x"0920";
    tmp(38481) := x"0920";
    tmp(38482) := x"0920";
    tmp(38483) := x"0920";
    tmp(38484) := x"0920";
    tmp(38485) := x"0900";
    tmp(38486) := x"0900";
    tmp(38487) := x"0900";
    tmp(38488) := x"08e0";
    tmp(38489) := x"0900";
    tmp(38490) := x"0900";
    tmp(38491) := x"0900";
    tmp(38492) := x"0900";
    tmp(38493) := x"1121";
    tmp(38494) := x"1141";
    tmp(38495) := x"1141";
    tmp(38496) := x"1141";
    tmp(38497) := x"1141";
    tmp(38498) := x"1121";
    tmp(38499) := x"0920";
    tmp(38500) := x"0920";
    tmp(38501) := x"0900";
    tmp(38502) := x"0920";
    tmp(38503) := x"0900";
    tmp(38504) := x"0900";
    tmp(38505) := x"0900";
    tmp(38506) := x"08e0";
    tmp(38507) := x"08e0";
    tmp(38508) := x"08e0";
    tmp(38509) := x"08e0";
    tmp(38510) := x"08e0";
    tmp(38511) := x"08e0";
    tmp(38512) := x"08e0";
    tmp(38513) := x"08e0";
    tmp(38514) := x"08e0";
    tmp(38515) := x"08e0";
    tmp(38516) := x"08e0";
    tmp(38517) := x"08c0";
    tmp(38518) := x"08c0";
    tmp(38519) := x"08c0";
    tmp(38520) := x"08c0";
    tmp(38521) := x"08e0";
    tmp(38522) := x"08e0";
    tmp(38523) := x"08c0";
    tmp(38524) := x"08c0";
    tmp(38525) := x"08c0";
    tmp(38526) := x"08a0";
    tmp(38527) := x"08c0";
    tmp(38528) := x"08c0";
    tmp(38529) := x"08c0";
    tmp(38530) := x"08c0";
    tmp(38531) := x"08c0";
    tmp(38532) := x"08c0";
    tmp(38533) := x"08e0";
    tmp(38534) := x"0900";
    tmp(38535) := x"0900";
    tmp(38536) := x"0900";
    tmp(38537) := x"0900";
    tmp(38538) := x"08e0";
    tmp(38539) := x"08e0";
    tmp(38540) := x"08e0";
    tmp(38541) := x"08c0";
    tmp(38542) := x"08c0";
    tmp(38543) := x"08c0";
    tmp(38544) := x"08c0";
    tmp(38545) := x"08c0";
    tmp(38546) := x"08a0";
    tmp(38547) := x"08a0";
    tmp(38548) := x"10a0";
    tmp(38549) := x"1080";
    tmp(38550) := x"1080";
    tmp(38551) := x"1080";
    tmp(38552) := x"1060";
    tmp(38553) := x"1060";
    tmp(38554) := x"1060";
    tmp(38555) := x"1060";
    tmp(38556) := x"1060";
    tmp(38557) := x"1060";
    tmp(38558) := x"1060";
    tmp(38559) := x"1060";
    tmp(38560) := x"1060";
    tmp(38561) := x"1060";
    tmp(38562) := x"1060";
    tmp(38563) := x"1060";
    tmp(38564) := x"1060";
    tmp(38565) := x"1060";
    tmp(38566) := x"1060";
    tmp(38567) := x"1060";
    tmp(38568) := x"1060";
    tmp(38569) := x"1040";
    tmp(38570) := x"1040";
    tmp(38571) := x"1040";
    tmp(38572) := x"1040";
    tmp(38573) := x"1040";
    tmp(38574) := x"1060";
    tmp(38575) := x"1060";
    tmp(38576) := x"1060";
    tmp(38577) := x"1060";
    tmp(38578) := x"1061";
    tmp(38579) := x"1061";
    tmp(38580) := x"1060";
    tmp(38581) := x"1061";
    tmp(38582) := x"1061";
    tmp(38583) := x"1061";
    tmp(38584) := x"1061";
    tmp(38585) := x"1061";
    tmp(38586) := x"1061";
    tmp(38587) := x"1061";
    tmp(38588) := x"1061";
    tmp(38589) := x"1060";
    tmp(38590) := x"1060";
    tmp(38591) := x"1040";
    tmp(38592) := x"1040";
    tmp(38593) := x"1040";
    tmp(38594) := x"1040";
    tmp(38595) := x"1040";
    tmp(38596) := x"1040";
    tmp(38597) := x"07e0";
    tmp(38598) := x"07e0";
    tmp(38599) := x"07e0";
    tmp(38600) := x"07e0";
    tmp(38601) := x"07e0";
    tmp(38602) := x"07e0";
    tmp(38603) := x"07e0";
    tmp(38604) := x"07e0";
    tmp(38605) := x"07e0";
    tmp(38606) := x"07e0";
    tmp(38607) := x"07e0";
    tmp(38608) := x"07e0";
    tmp(38609) := x"07e0";
    tmp(38610) := x"07e0";
    tmp(38611) := x"07e0";
    tmp(38612) := x"07e0";
    tmp(38613) := x"07e0";
    tmp(38614) := x"07e0";
    tmp(38615) := x"07e0";
    tmp(38616) := x"07e0";
    tmp(38617) := x"07e0";
    tmp(38618) := x"07e0";
    tmp(38619) := x"07e0";
    tmp(38620) := x"07e0";
    tmp(38621) := x"07e0";
    tmp(38622) := x"07e0";
    tmp(38623) := x"07e0";
    tmp(38624) := x"07e0";
    tmp(38625) := x"07e0";
    tmp(38626) := x"07e0";
    tmp(38627) := x"07e0";
    tmp(38628) := x"07e0";
    tmp(38629) := x"07e0";
    tmp(38630) := x"07e0";
    tmp(38631) := x"07e0";
    tmp(38632) := x"07e0";
    tmp(38633) := x"07e0";
    tmp(38634) := x"07e0";
    tmp(38635) := x"07e0";
    tmp(38636) := x"07e0";
    tmp(38637) := x"1060";
    tmp(38638) := x"1061";
    tmp(38639) := x"1061";
    tmp(38640) := x"0021";
    tmp(38641) := x"0a0a";
    tmp(38642) := x"0a09";
    tmp(38643) := x"0987";
    tmp(38644) := x"00c4";
    tmp(38645) := x"0061";
    tmp(38646) := x"0061";
    tmp(38647) := x"00a2";
    tmp(38648) := x"08a2";
    tmp(38649) := x"0082";
    tmp(38650) := x"0061";
    tmp(38651) := x"0021";
    tmp(38652) := x"0020";
    tmp(38653) := x"0000";
    tmp(38654) := x"0000";
    tmp(38655) := x"0000";
    tmp(38656) := x"0020";
    tmp(38657) := x"0860";
    tmp(38658) := x"08e1";
    tmp(38659) := x"1141";
    tmp(38660) := x"1141";
    tmp(38661) := x"1161";
    tmp(38662) := x"1161";
    tmp(38663) := x"1140";
    tmp(38664) := x"1120";
    tmp(38665) := x"1120";
    tmp(38666) := x"1120";
    tmp(38667) := x"1140";
    tmp(38668) := x"1120";
    tmp(38669) := x"1120";
    tmp(38670) := x"1140";
    tmp(38671) := x"1140";
    tmp(38672) := x"1140";
    tmp(38673) := x"1140";
    tmp(38674) := x"1141";
    tmp(38675) := x"1141";
    tmp(38676) := x"1141";
    tmp(38677) := x"1141";
    tmp(38678) := x"1161";
    tmp(38679) := x"1161";
    tmp(38680) := x"1161";
    tmp(38681) := x"1181";
    tmp(38682) := x"1181";
    tmp(38683) := x"1981";
    tmp(38684) := x"1981";
    tmp(38685) := x"1181";
    tmp(38686) := x"1181";
    tmp(38687) := x"1161";
    tmp(38688) := x"1161";
    tmp(38689) := x"1181";
    tmp(38690) := x"1161";
    tmp(38691) := x"1161";
    tmp(38692) := x"1181";
    tmp(38693) := x"1161";
    tmp(38694) := x"1161";
    tmp(38695) := x"1161";
    tmp(38696) := x"1161";
    tmp(38697) := x"1161";
    tmp(38698) := x"1141";
    tmp(38699) := x"1161";
    tmp(38700) := x"1161";
    tmp(38701) := x"1141";
    tmp(38702) := x"1161";
    tmp(38703) := x"1161";
    tmp(38704) := x"1161";
    tmp(38705) := x"1140";
    tmp(38706) := x"1140";
    tmp(38707) := x"1141";
    tmp(38708) := x"1141";
    tmp(38709) := x"1141";
    tmp(38710) := x"1141";
    tmp(38711) := x"1141";
    tmp(38712) := x"1161";
    tmp(38713) := x"1161";
    tmp(38714) := x"1141";
    tmp(38715) := x"1141";
    tmp(38716) := x"1140";
    tmp(38717) := x"1140";
    tmp(38718) := x"1140";
    tmp(38719) := x"1140";
    tmp(38720) := x"0920";
    tmp(38721) := x"0920";
    tmp(38722) := x"0920";
    tmp(38723) := x"0920";
    tmp(38724) := x"0920";
    tmp(38725) := x"0900";
    tmp(38726) := x"0900";
    tmp(38727) := x"0900";
    tmp(38728) := x"08e0";
    tmp(38729) := x"08e0";
    tmp(38730) := x"0900";
    tmp(38731) := x"0900";
    tmp(38732) := x"0920";
    tmp(38733) := x"1140";
    tmp(38734) := x"1141";
    tmp(38735) := x"1141";
    tmp(38736) := x"1141";
    tmp(38737) := x"1141";
    tmp(38738) := x"0920";
    tmp(38739) := x"0920";
    tmp(38740) := x"0920";
    tmp(38741) := x"0920";
    tmp(38742) := x"0920";
    tmp(38743) := x"0900";
    tmp(38744) := x"0900";
    tmp(38745) := x"0900";
    tmp(38746) := x"08e0";
    tmp(38747) := x"08e0";
    tmp(38748) := x"08e0";
    tmp(38749) := x"08e0";
    tmp(38750) := x"08e0";
    tmp(38751) := x"08e0";
    tmp(38752) := x"08e0";
    tmp(38753) := x"08e0";
    tmp(38754) := x"08e0";
    tmp(38755) := x"08e0";
    tmp(38756) := x"08c0";
    tmp(38757) := x"08c0";
    tmp(38758) := x"08c0";
    tmp(38759) := x"08c0";
    tmp(38760) := x"08c0";
    tmp(38761) := x"08e0";
    tmp(38762) := x"08c0";
    tmp(38763) := x"08c0";
    tmp(38764) := x"08a0";
    tmp(38765) := x"08a0";
    tmp(38766) := x"08a0";
    tmp(38767) := x"08a0";
    tmp(38768) := x"08c0";
    tmp(38769) := x"08c0";
    tmp(38770) := x"08c0";
    tmp(38771) := x"08c0";
    tmp(38772) := x"08e0";
    tmp(38773) := x"08e0";
    tmp(38774) := x"08e0";
    tmp(38775) := x"0900";
    tmp(38776) := x"0900";
    tmp(38777) := x"0900";
    tmp(38778) := x"08e0";
    tmp(38779) := x"08e0";
    tmp(38780) := x"08c0";
    tmp(38781) := x"08e0";
    tmp(38782) := x"08c0";
    tmp(38783) := x"08c0";
    tmp(38784) := x"08c0";
    tmp(38785) := x"08a0";
    tmp(38786) := x"08a0";
    tmp(38787) := x"08a0";
    tmp(38788) := x"10a0";
    tmp(38789) := x"0880";
    tmp(38790) := x"1080";
    tmp(38791) := x"1060";
    tmp(38792) := x"1060";
    tmp(38793) := x"1060";
    tmp(38794) := x"1060";
    tmp(38795) := x"1060";
    tmp(38796) := x"1060";
    tmp(38797) := x"1060";
    tmp(38798) := x"1060";
    tmp(38799) := x"1060";
    tmp(38800) := x"1060";
    tmp(38801) := x"1060";
    tmp(38802) := x"1060";
    tmp(38803) := x"1060";
    tmp(38804) := x"1060";
    tmp(38805) := x"1060";
    tmp(38806) := x"1060";
    tmp(38807) := x"1060";
    tmp(38808) := x"1040";
    tmp(38809) := x"1040";
    tmp(38810) := x"1040";
    tmp(38811) := x"1040";
    tmp(38812) := x"1040";
    tmp(38813) := x"1040";
    tmp(38814) := x"1040";
    tmp(38815) := x"1060";
    tmp(38816) := x"1060";
    tmp(38817) := x"1060";
    tmp(38818) := x"1060";
    tmp(38819) := x"1061";
    tmp(38820) := x"1060";
    tmp(38821) := x"1060";
    tmp(38822) := x"1061";
    tmp(38823) := x"1061";
    tmp(38824) := x"1061";
    tmp(38825) := x"1061";
    tmp(38826) := x"1061";
    tmp(38827) := x"1061";
    tmp(38828) := x"1061";
    tmp(38829) := x"1061";
    tmp(38830) := x"1060";
    tmp(38831) := x"1060";
    tmp(38832) := x"1040";
    tmp(38833) := x"1040";
    tmp(38834) := x"1040";
    tmp(38835) := x"1040";
    tmp(38836) := x"0840";
    tmp(38837) := x"07e0";
    tmp(38838) := x"07e0";
    tmp(38839) := x"07e0";
    tmp(38840) := x"07e0";
    tmp(38841) := x"07e0";
    tmp(38842) := x"07e0";
    tmp(38843) := x"07e0";
    tmp(38844) := x"07e0";
    tmp(38845) := x"07e0";
    tmp(38846) := x"07e0";
    tmp(38847) := x"07e0";
    tmp(38848) := x"07e0";
    tmp(38849) := x"07e0";
    tmp(38850) := x"07e0";
    tmp(38851) := x"07e0";
    tmp(38852) := x"07e0";
    tmp(38853) := x"07e0";
    tmp(38854) := x"07e0";
    tmp(38855) := x"07e0";
    tmp(38856) := x"07e0";
    tmp(38857) := x"07e0";
    tmp(38858) := x"07e0";
    tmp(38859) := x"07e0";
    tmp(38860) := x"07e0";
    tmp(38861) := x"07e0";
    tmp(38862) := x"07e0";
    tmp(38863) := x"07e0";
    tmp(38864) := x"07e0";
    tmp(38865) := x"07e0";
    tmp(38866) := x"07e0";
    tmp(38867) := x"07e0";
    tmp(38868) := x"07e0";
    tmp(38869) := x"07e0";
    tmp(38870) := x"07e0";
    tmp(38871) := x"07e0";
    tmp(38872) := x"07e0";
    tmp(38873) := x"07e0";
    tmp(38874) := x"07e0";
    tmp(38875) := x"07e0";
    tmp(38876) := x"07e0";
    tmp(38877) := x"1060";
    tmp(38878) := x"1061";
    tmp(38879) := x"1060";
    tmp(38880) := x"0020";
    tmp(38881) := x"00c3";
    tmp(38882) := x"0062";
    tmp(38883) := x"0061";
    tmp(38884) := x"0061";
    tmp(38885) := x"0082";
    tmp(38886) := x"0062";
    tmp(38887) := x"0041";
    tmp(38888) := x"0020";
    tmp(38889) := x"0000";
    tmp(38890) := x"0000";
    tmp(38891) := x"0000";
    tmp(38892) := x"0000";
    tmp(38893) := x"0000";
    tmp(38894) := x"0020";
    tmp(38895) := x"0040";
    tmp(38896) := x"08a0";
    tmp(38897) := x"08e0";
    tmp(38898) := x"0920";
    tmp(38899) := x"1120";
    tmp(38900) := x"1140";
    tmp(38901) := x"1140";
    tmp(38902) := x"1140";
    tmp(38903) := x"1140";
    tmp(38904) := x"1120";
    tmp(38905) := x"1120";
    tmp(38906) := x"1120";
    tmp(38907) := x"1120";
    tmp(38908) := x"1120";
    tmp(38909) := x"1120";
    tmp(38910) := x"1120";
    tmp(38911) := x"1120";
    tmp(38912) := x"1120";
    tmp(38913) := x"1120";
    tmp(38914) := x"1141";
    tmp(38915) := x"1141";
    tmp(38916) := x"1141";
    tmp(38917) := x"1141";
    tmp(38918) := x"1161";
    tmp(38919) := x"1161";
    tmp(38920) := x"1161";
    tmp(38921) := x"1161";
    tmp(38922) := x"1981";
    tmp(38923) := x"1181";
    tmp(38924) := x"1981";
    tmp(38925) := x"1181";
    tmp(38926) := x"1161";
    tmp(38927) := x"1181";
    tmp(38928) := x"1181";
    tmp(38929) := x"1181";
    tmp(38930) := x"1161";
    tmp(38931) := x"1161";
    tmp(38932) := x"1161";
    tmp(38933) := x"1161";
    tmp(38934) := x"1161";
    tmp(38935) := x"1161";
    tmp(38936) := x"1161";
    tmp(38937) := x"1161";
    tmp(38938) := x"1161";
    tmp(38939) := x"1161";
    tmp(38940) := x"1161";
    tmp(38941) := x"1161";
    tmp(38942) := x"1161";
    tmp(38943) := x"1161";
    tmp(38944) := x"1161";
    tmp(38945) := x"1161";
    tmp(38946) := x"1140";
    tmp(38947) := x"1140";
    tmp(38948) := x"1140";
    tmp(38949) := x"1141";
    tmp(38950) := x"1160";
    tmp(38951) := x"1161";
    tmp(38952) := x"1141";
    tmp(38953) := x"1161";
    tmp(38954) := x"1161";
    tmp(38955) := x"1141";
    tmp(38956) := x"1141";
    tmp(38957) := x"1140";
    tmp(38958) := x"1160";
    tmp(38959) := x"1140";
    tmp(38960) := x"1140";
    tmp(38961) := x"0920";
    tmp(38962) := x"0920";
    tmp(38963) := x"0920";
    tmp(38964) := x"0920";
    tmp(38965) := x"0900";
    tmp(38966) := x"0900";
    tmp(38967) := x"0900";
    tmp(38968) := x"0900";
    tmp(38969) := x"0900";
    tmp(38970) := x"08e0";
    tmp(38971) := x"0900";
    tmp(38972) := x"0920";
    tmp(38973) := x"0920";
    tmp(38974) := x"1140";
    tmp(38975) := x"1140";
    tmp(38976) := x"1140";
    tmp(38977) := x"0940";
    tmp(38978) := x"0940";
    tmp(38979) := x"0920";
    tmp(38980) := x"0920";
    tmp(38981) := x"0920";
    tmp(38982) := x"0900";
    tmp(38983) := x"0900";
    tmp(38984) := x"0900";
    tmp(38985) := x"0900";
    tmp(38986) := x"08e0";
    tmp(38987) := x"08e0";
    tmp(38988) := x"08e0";
    tmp(38989) := x"08e0";
    tmp(38990) := x"08e0";
    tmp(38991) := x"08e0";
    tmp(38992) := x"08e0";
    tmp(38993) := x"08e0";
    tmp(38994) := x"08e0";
    tmp(38995) := x"08e0";
    tmp(38996) := x"08e0";
    tmp(38997) := x"08c0";
    tmp(38998) := x"08c0";
    tmp(38999) := x"08c0";
    tmp(39000) := x"08c0";
    tmp(39001) := x"08c0";
    tmp(39002) := x"08c0";
    tmp(39003) := x"08c0";
    tmp(39004) := x"08c0";
    tmp(39005) := x"08a0";
    tmp(39006) := x"08a0";
    tmp(39007) := x"08c0";
    tmp(39008) := x"08a0";
    tmp(39009) := x"08c0";
    tmp(39010) := x"08c0";
    tmp(39011) := x"08c0";
    tmp(39012) := x"08c0";
    tmp(39013) := x"08c0";
    tmp(39014) := x"08e0";
    tmp(39015) := x"0900";
    tmp(39016) := x"0900";
    tmp(39017) := x"08e0";
    tmp(39018) := x"08e0";
    tmp(39019) := x"08e0";
    tmp(39020) := x"08e0";
    tmp(39021) := x"08c0";
    tmp(39022) := x"08c0";
    tmp(39023) := x"08c0";
    tmp(39024) := x"08c0";
    tmp(39025) := x"08c0";
    tmp(39026) := x"08a0";
    tmp(39027) := x"08a0";
    tmp(39028) := x"10a0";
    tmp(39029) := x"1080";
    tmp(39030) := x"1080";
    tmp(39031) := x"1080";
    tmp(39032) := x"1060";
    tmp(39033) := x"1060";
    tmp(39034) := x"1060";
    tmp(39035) := x"1060";
    tmp(39036) := x"1060";
    tmp(39037) := x"1060";
    tmp(39038) := x"1060";
    tmp(39039) := x"1060";
    tmp(39040) := x"1060";
    tmp(39041) := x"1060";
    tmp(39042) := x"1060";
    tmp(39043) := x"1060";
    tmp(39044) := x"1060";
    tmp(39045) := x"1060";
    tmp(39046) := x"1060";
    tmp(39047) := x"1040";
    tmp(39048) := x"1040";
    tmp(39049) := x"1040";
    tmp(39050) := x"1040";
    tmp(39051) := x"1040";
    tmp(39052) := x"1040";
    tmp(39053) := x"1040";
    tmp(39054) := x"1040";
    tmp(39055) := x"1060";
    tmp(39056) := x"1060";
    tmp(39057) := x"1060";
    tmp(39058) := x"1060";
    tmp(39059) := x"1061";
    tmp(39060) := x"1060";
    tmp(39061) := x"1061";
    tmp(39062) := x"1061";
    tmp(39063) := x"1061";
    tmp(39064) := x"1061";
    tmp(39065) := x"1061";
    tmp(39066) := x"1061";
    tmp(39067) := x"1061";
    tmp(39068) := x"1060";
    tmp(39069) := x"1060";
    tmp(39070) := x"1060";
    tmp(39071) := x"1060";
    tmp(39072) := x"1040";
    tmp(39073) := x"1040";
    tmp(39074) := x"0840";
    tmp(39075) := x"1040";
    tmp(39076) := x"0840";
    tmp(39077) := x"07e0";
    tmp(39078) := x"07e0";
    tmp(39079) := x"07e0";
    tmp(39080) := x"07e0";
    tmp(39081) := x"07e0";
    tmp(39082) := x"07e0";
    tmp(39083) := x"07e0";
    tmp(39084) := x"07e0";
    tmp(39085) := x"07e0";
    tmp(39086) := x"07e0";
    tmp(39087) := x"07e0";
    tmp(39088) := x"07e0";
    tmp(39089) := x"07e0";
    tmp(39090) := x"07e0";
    tmp(39091) := x"07e0";
    tmp(39092) := x"07e0";
    tmp(39093) := x"07e0";
    tmp(39094) := x"07e0";
    tmp(39095) := x"07e0";
    tmp(39096) := x"07e0";
    tmp(39097) := x"07e0";
    tmp(39098) := x"07e0";
    tmp(39099) := x"07e0";
    tmp(39100) := x"07e0";
    tmp(39101) := x"07e0";
    tmp(39102) := x"07e0";
    tmp(39103) := x"07e0";
    tmp(39104) := x"07e0";
    tmp(39105) := x"07e0";
    tmp(39106) := x"07e0";
    tmp(39107) := x"07e0";
    tmp(39108) := x"07e0";
    tmp(39109) := x"07e0";
    tmp(39110) := x"07e0";
    tmp(39111) := x"07e0";
    tmp(39112) := x"07e0";
    tmp(39113) := x"07e0";
    tmp(39114) := x"07e0";
    tmp(39115) := x"07e0";
    tmp(39116) := x"07e0";
    tmp(39117) := x"1061";
    tmp(39118) := x"1060";
    tmp(39119) := x"1061";
    tmp(39120) := x"0000";
    tmp(39121) := x"0020";
    tmp(39122) := x"0020";
    tmp(39123) := x"0020";
    tmp(39124) := x"0000";
    tmp(39125) := x"0000";
    tmp(39126) := x"0000";
    tmp(39127) := x"0000";
    tmp(39128) := x"0000";
    tmp(39129) := x"0000";
    tmp(39130) := x"0000";
    tmp(39131) := x"0000";
    tmp(39132) := x"0020";
    tmp(39133) := x"0040";
    tmp(39134) := x"0880";
    tmp(39135) := x"08c0";
    tmp(39136) := x"08e0";
    tmp(39137) := x"08e0";
    tmp(39138) := x"0900";
    tmp(39139) := x"0920";
    tmp(39140) := x"1120";
    tmp(39141) := x"1120";
    tmp(39142) := x"1120";
    tmp(39143) := x"1120";
    tmp(39144) := x"1120";
    tmp(39145) := x"0920";
    tmp(39146) := x"0900";
    tmp(39147) := x"0900";
    tmp(39148) := x"0920";
    tmp(39149) := x"1120";
    tmp(39150) := x"1120";
    tmp(39151) := x"1120";
    tmp(39152) := x"1120";
    tmp(39153) := x"1140";
    tmp(39154) := x"1140";
    tmp(39155) := x"1141";
    tmp(39156) := x"1141";
    tmp(39157) := x"1141";
    tmp(39158) := x"1141";
    tmp(39159) := x"1161";
    tmp(39160) := x"1161";
    tmp(39161) := x"1161";
    tmp(39162) := x"1181";
    tmp(39163) := x"1981";
    tmp(39164) := x"1181";
    tmp(39165) := x"1181";
    tmp(39166) := x"1161";
    tmp(39167) := x"1161";
    tmp(39168) := x"1161";
    tmp(39169) := x"1181";
    tmp(39170) := x"1181";
    tmp(39171) := x"1161";
    tmp(39172) := x"1161";
    tmp(39173) := x"1161";
    tmp(39174) := x"1161";
    tmp(39175) := x"1161";
    tmp(39176) := x"1161";
    tmp(39177) := x"1161";
    tmp(39178) := x"1161";
    tmp(39179) := x"1161";
    tmp(39180) := x"1161";
    tmp(39181) := x"1161";
    tmp(39182) := x"1161";
    tmp(39183) := x"1161";
    tmp(39184) := x"1161";
    tmp(39185) := x"1140";
    tmp(39186) := x"1140";
    tmp(39187) := x"1140";
    tmp(39188) := x"1140";
    tmp(39189) := x"1140";
    tmp(39190) := x"1161";
    tmp(39191) := x"1141";
    tmp(39192) := x"1161";
    tmp(39193) := x"1161";
    tmp(39194) := x"1161";
    tmp(39195) := x"1161";
    tmp(39196) := x"1141";
    tmp(39197) := x"1161";
    tmp(39198) := x"1160";
    tmp(39199) := x"1140";
    tmp(39200) := x"1140";
    tmp(39201) := x"1140";
    tmp(39202) := x"0920";
    tmp(39203) := x"0920";
    tmp(39204) := x"0920";
    tmp(39205) := x"0900";
    tmp(39206) := x"0900";
    tmp(39207) := x"0900";
    tmp(39208) := x"0900";
    tmp(39209) := x"08e0";
    tmp(39210) := x"08e0";
    tmp(39211) := x"08e0";
    tmp(39212) := x"08e0";
    tmp(39213) := x"0900";
    tmp(39214) := x"0920";
    tmp(39215) := x"0920";
    tmp(39216) := x"0920";
    tmp(39217) := x"0900";
    tmp(39218) := x"0920";
    tmp(39219) := x"0920";
    tmp(39220) := x"0900";
    tmp(39221) := x"0900";
    tmp(39222) := x"0900";
    tmp(39223) := x"0900";
    tmp(39224) := x"0900";
    tmp(39225) := x"08e0";
    tmp(39226) := x"0900";
    tmp(39227) := x"0900";
    tmp(39228) := x"0900";
    tmp(39229) := x"08e0";
    tmp(39230) := x"08e0";
    tmp(39231) := x"08e0";
    tmp(39232) := x"08e0";
    tmp(39233) := x"08e0";
    tmp(39234) := x"08e0";
    tmp(39235) := x"08e0";
    tmp(39236) := x"08c0";
    tmp(39237) := x"08e0";
    tmp(39238) := x"08c0";
    tmp(39239) := x"08c0";
    tmp(39240) := x"08c0";
    tmp(39241) := x"08c0";
    tmp(39242) := x"08c0";
    tmp(39243) := x"08c0";
    tmp(39244) := x"08c0";
    tmp(39245) := x"08a0";
    tmp(39246) := x"08a0";
    tmp(39247) := x"08a0";
    tmp(39248) := x"08a0";
    tmp(39249) := x"08c0";
    tmp(39250) := x"08c0";
    tmp(39251) := x"08c0";
    tmp(39252) := x"08c0";
    tmp(39253) := x"08c0";
    tmp(39254) := x"08e0";
    tmp(39255) := x"08e0";
    tmp(39256) := x"08e0";
    tmp(39257) := x"08e0";
    tmp(39258) := x"08e0";
    tmp(39259) := x"08e0";
    tmp(39260) := x"08e0";
    tmp(39261) := x"08e0";
    tmp(39262) := x"08c0";
    tmp(39263) := x"08c0";
    tmp(39264) := x"08c0";
    tmp(39265) := x"08c0";
    tmp(39266) := x"08a0";
    tmp(39267) := x"08a0";
    tmp(39268) := x"08a0";
    tmp(39269) := x"1080";
    tmp(39270) := x"1080";
    tmp(39271) := x"1060";
    tmp(39272) := x"1060";
    tmp(39273) := x"1060";
    tmp(39274) := x"1060";
    tmp(39275) := x"1060";
    tmp(39276) := x"1060";
    tmp(39277) := x"1060";
    tmp(39278) := x"1060";
    tmp(39279) := x"1060";
    tmp(39280) := x"1060";
    tmp(39281) := x"1060";
    tmp(39282) := x"1060";
    tmp(39283) := x"1060";
    tmp(39284) := x"1060";
    tmp(39285) := x"1060";
    tmp(39286) := x"1060";
    tmp(39287) := x"1040";
    tmp(39288) := x"1040";
    tmp(39289) := x"1040";
    tmp(39290) := x"1040";
    tmp(39291) := x"1040";
    tmp(39292) := x"1040";
    tmp(39293) := x"1060";
    tmp(39294) := x"1040";
    tmp(39295) := x"1060";
    tmp(39296) := x"1060";
    tmp(39297) := x"1061";
    tmp(39298) := x"1061";
    tmp(39299) := x"1060";
    tmp(39300) := x"1061";
    tmp(39301) := x"1061";
    tmp(39302) := x"1061";
    tmp(39303) := x"1061";
    tmp(39304) := x"1061";
    tmp(39305) := x"1061";
    tmp(39306) := x"1061";
    tmp(39307) := x"1061";
    tmp(39308) := x"1061";
    tmp(39309) := x"1060";
    tmp(39310) := x"1060";
    tmp(39311) := x"1040";
    tmp(39312) := x"1040";
    tmp(39313) := x"1040";
    tmp(39314) := x"1040";
    tmp(39315) := x"1040";
    tmp(39316) := x"0840";
    tmp(39317) := x"07e0";
    tmp(39318) := x"07e0";
    tmp(39319) := x"07e0";
    tmp(39320) := x"07e0";
    tmp(39321) := x"07e0";
    tmp(39322) := x"07e0";
    tmp(39323) := x"07e0";
    tmp(39324) := x"07e0";
    tmp(39325) := x"07e0";
    tmp(39326) := x"07e0";
    tmp(39327) := x"07e0";
    tmp(39328) := x"07e0";
    tmp(39329) := x"07e0";
    tmp(39330) := x"07e0";
    tmp(39331) := x"07e0";
    tmp(39332) := x"07e0";
    tmp(39333) := x"07e0";
    tmp(39334) := x"07e0";
    tmp(39335) := x"07e0";
    tmp(39336) := x"07e0";
    tmp(39337) := x"07e0";
    tmp(39338) := x"07e0";
    tmp(39339) := x"07e0";
    tmp(39340) := x"07e0";
    tmp(39341) := x"07e0";
    tmp(39342) := x"07e0";
    tmp(39343) := x"07e0";
    tmp(39344) := x"07e0";
    tmp(39345) := x"07e0";
    tmp(39346) := x"07e0";
    tmp(39347) := x"07e0";
    tmp(39348) := x"07e0";
    tmp(39349) := x"07e0";
    tmp(39350) := x"07e0";
    tmp(39351) := x"07e0";
    tmp(39352) := x"07e0";
    tmp(39353) := x"07e0";
    tmp(39354) := x"07e0";
    tmp(39355) := x"07e0";
    tmp(39356) := x"07e0";
    tmp(39357) := x"1061";
    tmp(39358) := x"1061";
    tmp(39359) := x"1061";
    tmp(39360) := x"0000";
    tmp(39361) := x"0000";
    tmp(39362) := x"0000";
    tmp(39363) := x"0000";
    tmp(39364) := x"0000";
    tmp(39365) := x"0000";
    tmp(39366) := x"0000";
    tmp(39367) := x"0000";
    tmp(39368) := x"0000";
    tmp(39369) := x"0000";
    tmp(39370) := x"0020";
    tmp(39371) := x"0040";
    tmp(39372) := x"0860";
    tmp(39373) := x"08a0";
    tmp(39374) := x"08c0";
    tmp(39375) := x"08c0";
    tmp(39376) := x"08c0";
    tmp(39377) := x"08c0";
    tmp(39378) := x"08e0";
    tmp(39379) := x"0900";
    tmp(39380) := x"0900";
    tmp(39381) := x"0920";
    tmp(39382) := x"0920";
    tmp(39383) := x"0920";
    tmp(39384) := x"0920";
    tmp(39385) := x"0900";
    tmp(39386) := x"0900";
    tmp(39387) := x"0920";
    tmp(39388) := x"0900";
    tmp(39389) := x"0920";
    tmp(39390) := x"0920";
    tmp(39391) := x"0920";
    tmp(39392) := x"0920";
    tmp(39393) := x"1140";
    tmp(39394) := x"1140";
    tmp(39395) := x"1140";
    tmp(39396) := x"1141";
    tmp(39397) := x"1141";
    tmp(39398) := x"1141";
    tmp(39399) := x"1161";
    tmp(39400) := x"1161";
    tmp(39401) := x"1161";
    tmp(39402) := x"1181";
    tmp(39403) := x"1161";
    tmp(39404) := x"1161";
    tmp(39405) := x"1161";
    tmp(39406) := x"1161";
    tmp(39407) := x"1161";
    tmp(39408) := x"1161";
    tmp(39409) := x"1161";
    tmp(39410) := x"1181";
    tmp(39411) := x"1161";
    tmp(39412) := x"1161";
    tmp(39413) := x"1161";
    tmp(39414) := x"1161";
    tmp(39415) := x"1161";
    tmp(39416) := x"1161";
    tmp(39417) := x"1161";
    tmp(39418) := x"1181";
    tmp(39419) := x"1161";
    tmp(39420) := x"1161";
    tmp(39421) := x"1161";
    tmp(39422) := x"1161";
    tmp(39423) := x"1161";
    tmp(39424) := x"1161";
    tmp(39425) := x"1140";
    tmp(39426) := x"1140";
    tmp(39427) := x"1140";
    tmp(39428) := x"1140";
    tmp(39429) := x"1140";
    tmp(39430) := x"1141";
    tmp(39431) := x"1141";
    tmp(39432) := x"1161";
    tmp(39433) := x"1161";
    tmp(39434) := x"1181";
    tmp(39435) := x"1161";
    tmp(39436) := x"1161";
    tmp(39437) := x"1181";
    tmp(39438) := x"1160";
    tmp(39439) := x"1140";
    tmp(39440) := x"1140";
    tmp(39441) := x"0940";
    tmp(39442) := x"0920";
    tmp(39443) := x"0920";
    tmp(39444) := x"0920";
    tmp(39445) := x"0920";
    tmp(39446) := x"0900";
    tmp(39447) := x"0900";
    tmp(39448) := x"0900";
    tmp(39449) := x"0900";
    tmp(39450) := x"08e0";
    tmp(39451) := x"08e0";
    tmp(39452) := x"08e0";
    tmp(39453) := x"08e0";
    tmp(39454) := x"0900";
    tmp(39455) := x"0900";
    tmp(39456) := x"0900";
    tmp(39457) := x"0900";
    tmp(39458) := x"0900";
    tmp(39459) := x"0900";
    tmp(39460) := x"0900";
    tmp(39461) := x"0900";
    tmp(39462) := x"0900";
    tmp(39463) := x"0900";
    tmp(39464) := x"0900";
    tmp(39465) := x"0900";
    tmp(39466) := x"0900";
    tmp(39467) := x"08e0";
    tmp(39468) := x"08e0";
    tmp(39469) := x"08e0";
    tmp(39470) := x"08e0";
    tmp(39471) := x"08e0";
    tmp(39472) := x"08e0";
    tmp(39473) := x"08e0";
    tmp(39474) := x"08e0";
    tmp(39475) := x"08c0";
    tmp(39476) := x"08c0";
    tmp(39477) := x"08c0";
    tmp(39478) := x"08c0";
    tmp(39479) := x"08c0";
    tmp(39480) := x"08a0";
    tmp(39481) := x"08c0";
    tmp(39482) := x"08c0";
    tmp(39483) := x"08a0";
    tmp(39484) := x"08a0";
    tmp(39485) := x"08a0";
    tmp(39486) := x"08a0";
    tmp(39487) := x"08a0";
    tmp(39488) := x"08a0";
    tmp(39489) := x"08a0";
    tmp(39490) := x"08c0";
    tmp(39491) := x"08c0";
    tmp(39492) := x"08c0";
    tmp(39493) := x"08c0";
    tmp(39494) := x"08e0";
    tmp(39495) := x"08e0";
    tmp(39496) := x"08e0";
    tmp(39497) := x"08e0";
    tmp(39498) := x"08e0";
    tmp(39499) := x"08e0";
    tmp(39500) := x"08e0";
    tmp(39501) := x"08c0";
    tmp(39502) := x"08c0";
    tmp(39503) := x"08c0";
    tmp(39504) := x"08c0";
    tmp(39505) := x"08a0";
    tmp(39506) := x"08a0";
    tmp(39507) := x"08a0";
    tmp(39508) := x"0880";
    tmp(39509) := x"1080";
    tmp(39510) := x"0880";
    tmp(39511) := x"1080";
    tmp(39512) := x"1060";
    tmp(39513) := x"1060";
    tmp(39514) := x"1060";
    tmp(39515) := x"1060";
    tmp(39516) := x"1060";
    tmp(39517) := x"1060";
    tmp(39518) := x"1060";
    tmp(39519) := x"1060";
    tmp(39520) := x"1060";
    tmp(39521) := x"1060";
    tmp(39522) := x"1060";
    tmp(39523) := x"1060";
    tmp(39524) := x"1060";
    tmp(39525) := x"1060";
    tmp(39526) := x"1040";
    tmp(39527) := x"1040";
    tmp(39528) := x"1040";
    tmp(39529) := x"1040";
    tmp(39530) := x"1040";
    tmp(39531) := x"1040";
    tmp(39532) := x"1040";
    tmp(39533) := x"1060";
    tmp(39534) := x"1040";
    tmp(39535) := x"1060";
    tmp(39536) := x"1060";
    tmp(39537) := x"1060";
    tmp(39538) := x"1061";
    tmp(39539) := x"1060";
    tmp(39540) := x"1061";
    tmp(39541) := x"1061";
    tmp(39542) := x"1061";
    tmp(39543) := x"1061";
    tmp(39544) := x"1061";
    tmp(39545) := x"1061";
    tmp(39546) := x"1061";
    tmp(39547) := x"1061";
    tmp(39548) := x"1060";
    tmp(39549) := x"1061";
    tmp(39550) := x"1060";
    tmp(39551) := x"1040";
    tmp(39552) := x"1040";
    tmp(39553) := x"0840";
    tmp(39554) := x"0840";
    tmp(39555) := x"0840";
    tmp(39556) := x"0840";
    tmp(39557) := x"001f";
    tmp(39558) := x"001f";
    tmp(39559) := x"001f";
    tmp(39560) := x"001f";
    tmp(39561) := x"001f";
    tmp(39562) := x"001f";
    tmp(39563) := x"001f";
    tmp(39564) := x"001f";
    tmp(39565) := x"001f";
    tmp(39566) := x"001f";
    tmp(39567) := x"001f";
    tmp(39568) := x"001f";
    tmp(39569) := x"001f";
    tmp(39570) := x"001f";
    tmp(39571) := x"001f";
    tmp(39572) := x"001f";
    tmp(39573) := x"001f";
    tmp(39574) := x"001f";
    tmp(39575) := x"001f";
    tmp(39576) := x"001f";
    tmp(39577) := x"001f";
    tmp(39578) := x"001f";
    tmp(39579) := x"001f";
    tmp(39580) := x"001f";
    tmp(39581) := x"001f";
    tmp(39582) := x"001f";
    tmp(39583) := x"001f";
    tmp(39584) := x"001f";
    tmp(39585) := x"001f";
    tmp(39586) := x"001f";
    tmp(39587) := x"001f";
    tmp(39588) := x"001f";
    tmp(39589) := x"001f";
    tmp(39590) := x"001f";
    tmp(39591) := x"001f";
    tmp(39592) := x"001f";
    tmp(39593) := x"001f";
    tmp(39594) := x"001f";
    tmp(39595) := x"001f";
    tmp(39596) := x"001f";
    tmp(39597) := x"1061";
    tmp(39598) := x"1061";
    tmp(39599) := x"1061";
    tmp(39600) := x"0000";
    tmp(39601) := x"0000";
    tmp(39602) := x"0000";
    tmp(39603) := x"0000";
    tmp(39604) := x"0000";
    tmp(39605) := x"0000";
    tmp(39606) := x"0000";
    tmp(39607) := x"0020";
    tmp(39608) := x"0020";
    tmp(39609) := x"0040";
    tmp(39610) := x"0880";
    tmp(39611) := x"08a0";
    tmp(39612) := x"08a0";
    tmp(39613) := x"08a0";
    tmp(39614) := x"08c0";
    tmp(39615) := x"08c0";
    tmp(39616) := x"08c0";
    tmp(39617) := x"08c0";
    tmp(39618) := x"08c0";
    tmp(39619) := x"08e0";
    tmp(39620) := x"08e0";
    tmp(39621) := x"0900";
    tmp(39622) := x"0900";
    tmp(39623) := x"0900";
    tmp(39624) := x"0900";
    tmp(39625) := x"0900";
    tmp(39626) := x"0900";
    tmp(39627) := x"0900";
    tmp(39628) := x"0900";
    tmp(39629) := x"0920";
    tmp(39630) := x"0920";
    tmp(39631) := x"0920";
    tmp(39632) := x"0920";
    tmp(39633) := x"1120";
    tmp(39634) := x"1140";
    tmp(39635) := x"1140";
    tmp(39636) := x"1141";
    tmp(39637) := x"1141";
    tmp(39638) := x"1141";
    tmp(39639) := x"1141";
    tmp(39640) := x"1141";
    tmp(39641) := x"1161";
    tmp(39642) := x"1181";
    tmp(39643) := x"1181";
    tmp(39644) := x"1181";
    tmp(39645) := x"1161";
    tmp(39646) := x"1160";
    tmp(39647) := x"1161";
    tmp(39648) := x"1161";
    tmp(39649) := x"1161";
    tmp(39650) := x"1181";
    tmp(39651) := x"1181";
    tmp(39652) := x"1161";
    tmp(39653) := x"1161";
    tmp(39654) := x"1161";
    tmp(39655) := x"1161";
    tmp(39656) := x"1161";
    tmp(39657) := x"1161";
    tmp(39658) := x"1161";
    tmp(39659) := x"1160";
    tmp(39660) := x"1161";
    tmp(39661) := x"1161";
    tmp(39662) := x"1161";
    tmp(39663) := x"1161";
    tmp(39664) := x"1161";
    tmp(39665) := x"1140";
    tmp(39666) := x"0940";
    tmp(39667) := x"0920";
    tmp(39668) := x"1140";
    tmp(39669) := x"1140";
    tmp(39670) := x"1140";
    tmp(39671) := x"1160";
    tmp(39672) := x"1160";
    tmp(39673) := x"1161";
    tmp(39674) := x"1181";
    tmp(39675) := x"1161";
    tmp(39676) := x"1161";
    tmp(39677) := x"1160";
    tmp(39678) := x"1160";
    tmp(39679) := x"1160";
    tmp(39680) := x"1140";
    tmp(39681) := x"0940";
    tmp(39682) := x"0920";
    tmp(39683) := x"0920";
    tmp(39684) := x"0920";
    tmp(39685) := x"0900";
    tmp(39686) := x"0900";
    tmp(39687) := x"0900";
    tmp(39688) := x"0900";
    tmp(39689) := x"0900";
    tmp(39690) := x"08e0";
    tmp(39691) := x"08e0";
    tmp(39692) := x"08e0";
    tmp(39693) := x"08e0";
    tmp(39694) := x"0900";
    tmp(39695) := x"0900";
    tmp(39696) := x"0900";
    tmp(39697) := x"0900";
    tmp(39698) := x"0900";
    tmp(39699) := x"0900";
    tmp(39700) := x"0900";
    tmp(39701) := x"0900";
    tmp(39702) := x"0900";
    tmp(39703) := x"0900";
    tmp(39704) := x"0900";
    tmp(39705) := x"0900";
    tmp(39706) := x"08e0";
    tmp(39707) := x"08e0";
    tmp(39708) := x"08e0";
    tmp(39709) := x"08e0";
    tmp(39710) := x"08e0";
    tmp(39711) := x"08e0";
    tmp(39712) := x"08e0";
    tmp(39713) := x"08e0";
    tmp(39714) := x"08c0";
    tmp(39715) := x"08c0";
    tmp(39716) := x"08c0";
    tmp(39717) := x"08c0";
    tmp(39718) := x"08c0";
    tmp(39719) := x"08c0";
    tmp(39720) := x"08a0";
    tmp(39721) := x"08a0";
    tmp(39722) := x"08c0";
    tmp(39723) := x"08a0";
    tmp(39724) := x"08a0";
    tmp(39725) := x"08a0";
    tmp(39726) := x"08a0";
    tmp(39727) := x"08a0";
    tmp(39728) := x"08a0";
    tmp(39729) := x"08a0";
    tmp(39730) := x"08c0";
    tmp(39731) := x"08a0";
    tmp(39732) := x"08c0";
    tmp(39733) := x"08c0";
    tmp(39734) := x"08c0";
    tmp(39735) := x"08e0";
    tmp(39736) := x"08e0";
    tmp(39737) := x"08e0";
    tmp(39738) := x"08e0";
    tmp(39739) := x"08e0";
    tmp(39740) := x"08e0";
    tmp(39741) := x"08c0";
    tmp(39742) := x"08c0";
    tmp(39743) := x"08c0";
    tmp(39744) := x"08c0";
    tmp(39745) := x"08a0";
    tmp(39746) := x"08a0";
    tmp(39747) := x"08a0";
    tmp(39748) := x"10a0";
    tmp(39749) := x"0880";
    tmp(39750) := x"1080";
    tmp(39751) := x"1060";
    tmp(39752) := x"1060";
    tmp(39753) := x"1060";
    tmp(39754) := x"1060";
    tmp(39755) := x"0860";
    tmp(39756) := x"1060";
    tmp(39757) := x"1060";
    tmp(39758) := x"1060";
    tmp(39759) := x"1060";
    tmp(39760) := x"1060";
    tmp(39761) := x"1060";
    tmp(39762) := x"1060";
    tmp(39763) := x"1060";
    tmp(39764) := x"1060";
    tmp(39765) := x"1040";
    tmp(39766) := x"1040";
    tmp(39767) := x"1060";
    tmp(39768) := x"1040";
    tmp(39769) := x"1040";
    tmp(39770) := x"1040";
    tmp(39771) := x"1040";
    tmp(39772) := x"1060";
    tmp(39773) := x"1060";
    tmp(39774) := x"1040";
    tmp(39775) := x"1040";
    tmp(39776) := x"1060";
    tmp(39777) := x"1060";
    tmp(39778) := x"1060";
    tmp(39779) := x"1060";
    tmp(39780) := x"1061";
    tmp(39781) := x"1061";
    tmp(39782) := x"1061";
    tmp(39783) := x"1061";
    tmp(39784) := x"1061";
    tmp(39785) := x"1061";
    tmp(39786) := x"1061";
    tmp(39787) := x"1061";
    tmp(39788) := x"1061";
    tmp(39789) := x"1060";
    tmp(39790) := x"1040";
    tmp(39791) := x"1040";
    tmp(39792) := x"1040";
    tmp(39793) := x"0840";
    tmp(39794) := x"0840";
    tmp(39795) := x"0840";
    tmp(39796) := x"0840";
    tmp(39797) := x"001f";
    tmp(39798) := x"001f";
    tmp(39799) := x"001f";
    tmp(39800) := x"001f";
    tmp(39801) := x"001f";
    tmp(39802) := x"001f";
    tmp(39803) := x"001f";
    tmp(39804) := x"001f";
    tmp(39805) := x"001f";
    tmp(39806) := x"001f";
    tmp(39807) := x"001f";
    tmp(39808) := x"001f";
    tmp(39809) := x"001f";
    tmp(39810) := x"001f";
    tmp(39811) := x"001f";
    tmp(39812) := x"001f";
    tmp(39813) := x"001f";
    tmp(39814) := x"001f";
    tmp(39815) := x"001f";
    tmp(39816) := x"001f";
    tmp(39817) := x"001f";
    tmp(39818) := x"001f";
    tmp(39819) := x"001f";
    tmp(39820) := x"001f";
    tmp(39821) := x"001f";
    tmp(39822) := x"001f";
    tmp(39823) := x"001f";
    tmp(39824) := x"001f";
    tmp(39825) := x"001f";
    tmp(39826) := x"001f";
    tmp(39827) := x"001f";
    tmp(39828) := x"001f";
    tmp(39829) := x"001f";
    tmp(39830) := x"001f";
    tmp(39831) := x"001f";
    tmp(39832) := x"001f";
    tmp(39833) := x"001f";
    tmp(39834) := x"001f";
    tmp(39835) := x"001f";
    tmp(39836) := x"001f";
    tmp(39837) := x"1061";
    tmp(39838) := x"1061";
    tmp(39839) := x"1061";
    tmp(39840) := x"0000";
    tmp(39841) := x"0000";
    tmp(39842) := x"0000";
    tmp(39843) := x"0020";
    tmp(39844) := x"0020";
    tmp(39845) := x"0020";
    tmp(39846) := x"0020";
    tmp(39847) := x"0040";
    tmp(39848) := x"0860";
    tmp(39849) := x"0880";
    tmp(39850) := x"08a0";
    tmp(39851) := x"08a0";
    tmp(39852) := x"08a0";
    tmp(39853) := x"08a0";
    tmp(39854) := x"08a0";
    tmp(39855) := x"08c0";
    tmp(39856) := x"08c0";
    tmp(39857) := x"08c0";
    tmp(39858) := x"08c0";
    tmp(39859) := x"08c0";
    tmp(39860) := x"08e0";
    tmp(39861) := x"0900";
    tmp(39862) := x"0900";
    tmp(39863) := x"0900";
    tmp(39864) := x"0900";
    tmp(39865) := x"0900";
    tmp(39866) := x"0900";
    tmp(39867) := x"0900";
    tmp(39868) := x"0900";
    tmp(39869) := x"0920";
    tmp(39870) := x"0900";
    tmp(39871) := x"0900";
    tmp(39872) := x"0920";
    tmp(39873) := x"0920";
    tmp(39874) := x"1120";
    tmp(39875) := x"1140";
    tmp(39876) := x"1141";
    tmp(39877) := x"1141";
    tmp(39878) := x"1141";
    tmp(39879) := x"1141";
    tmp(39880) := x"1141";
    tmp(39881) := x"1161";
    tmp(39882) := x"1161";
    tmp(39883) := x"1181";
    tmp(39884) := x"1161";
    tmp(39885) := x"1161";
    tmp(39886) := x"1140";
    tmp(39887) := x"1140";
    tmp(39888) := x"1161";
    tmp(39889) := x"1161";
    tmp(39890) := x"1181";
    tmp(39891) := x"1161";
    tmp(39892) := x"1161";
    tmp(39893) := x"1161";
    tmp(39894) := x"1161";
    tmp(39895) := x"1161";
    tmp(39896) := x"1161";
    tmp(39897) := x"1161";
    tmp(39898) := x"1161";
    tmp(39899) := x"1161";
    tmp(39900) := x"1161";
    tmp(39901) := x"1141";
    tmp(39902) := x"1161";
    tmp(39903) := x"1161";
    tmp(39904) := x"1141";
    tmp(39905) := x"1140";
    tmp(39906) := x"1120";
    tmp(39907) := x"0920";
    tmp(39908) := x"0920";
    tmp(39909) := x"0920";
    tmp(39910) := x"0940";
    tmp(39911) := x"1140";
    tmp(39912) := x"1140";
    tmp(39913) := x"1140";
    tmp(39914) := x"1140";
    tmp(39915) := x"1140";
    tmp(39916) := x"1140";
    tmp(39917) := x"1140";
    tmp(39918) := x"1140";
    tmp(39919) := x"1140";
    tmp(39920) := x"1140";
    tmp(39921) := x"0920";
    tmp(39922) := x"0920";
    tmp(39923) := x"0920";
    tmp(39924) := x"0900";
    tmp(39925) := x"0900";
    tmp(39926) := x"0900";
    tmp(39927) := x"0900";
    tmp(39928) := x"0900";
    tmp(39929) := x"0900";
    tmp(39930) := x"08e0";
    tmp(39931) := x"0900";
    tmp(39932) := x"08e0";
    tmp(39933) := x"0900";
    tmp(39934) := x"08e0";
    tmp(39935) := x"0900";
    tmp(39936) := x"0900";
    tmp(39937) := x"0900";
    tmp(39938) := x"0900";
    tmp(39939) := x"0900";
    tmp(39940) := x"0900";
    tmp(39941) := x"0900";
    tmp(39942) := x"0900";
    tmp(39943) := x"0900";
    tmp(39944) := x"0900";
    tmp(39945) := x"0900";
    tmp(39946) := x"08e0";
    tmp(39947) := x"08e0";
    tmp(39948) := x"08e0";
    tmp(39949) := x"08e0";
    tmp(39950) := x"08e0";
    tmp(39951) := x"08e0";
    tmp(39952) := x"08e0";
    tmp(39953) := x"08e0";
    tmp(39954) := x"08e0";
    tmp(39955) := x"08c0";
    tmp(39956) := x"08c0";
    tmp(39957) := x"08c0";
    tmp(39958) := x"08c0";
    tmp(39959) := x"08c0";
    tmp(39960) := x"08a0";
    tmp(39961) := x"08a0";
    tmp(39962) := x"08c0";
    tmp(39963) := x"08a0";
    tmp(39964) := x"08a0";
    tmp(39965) := x"08a0";
    tmp(39966) := x"08a0";
    tmp(39967) := x"08a0";
    tmp(39968) := x"08a0";
    tmp(39969) := x"08a0";
    tmp(39970) := x"08a0";
    tmp(39971) := x"08a0";
    tmp(39972) := x"08a0";
    tmp(39973) := x"08c0";
    tmp(39974) := x"08c0";
    tmp(39975) := x"08e0";
    tmp(39976) := x"08e0";
    tmp(39977) := x"08c0";
    tmp(39978) := x"08e0";
    tmp(39979) := x"08c0";
    tmp(39980) := x"08c0";
    tmp(39981) := x"08c0";
    tmp(39982) := x"08c0";
    tmp(39983) := x"08c0";
    tmp(39984) := x"08a0";
    tmp(39985) := x"08a0";
    tmp(39986) := x"08a0";
    tmp(39987) := x"08a0";
    tmp(39988) := x"0880";
    tmp(39989) := x"0880";
    tmp(39990) := x"0880";
    tmp(39991) := x"1060";
    tmp(39992) := x"1060";
    tmp(39993) := x"1060";
    tmp(39994) := x"1060";
    tmp(39995) := x"1060";
    tmp(39996) := x"1060";
    tmp(39997) := x"1060";
    tmp(39998) := x"1060";
    tmp(39999) := x"1040";
    tmp(40000) := x"1860";
    tmp(40001) := x"1860";
    tmp(40002) := x"1040";
    tmp(40003) := x"1040";
    tmp(40004) := x"1040";
    tmp(40005) := x"1040";
    tmp(40006) := x"1040";
    tmp(40007) := x"1040";
    tmp(40008) := x"1040";
    tmp(40009) := x"1060";
    tmp(40010) := x"1040";
    tmp(40011) := x"1040";
    tmp(40012) := x"1060";
    tmp(40013) := x"1060";
    tmp(40014) := x"1040";
    tmp(40015) := x"1040";
    tmp(40016) := x"1040";
    tmp(40017) := x"1060";
    tmp(40018) := x"1060";
    tmp(40019) := x"1061";
    tmp(40020) := x"1061";
    tmp(40021) := x"1061";
    tmp(40022) := x"1061";
    tmp(40023) := x"1061";
    tmp(40024) := x"1061";
    tmp(40025) := x"1061";
    tmp(40026) := x"1061";
    tmp(40027) := x"1060";
    tmp(40028) := x"1060";
    tmp(40029) := x"1040";
    tmp(40030) := x"1040";
    tmp(40031) := x"0840";
    tmp(40032) := x"0840";
    tmp(40033) := x"0840";
    tmp(40034) := x"0840";
    tmp(40035) := x"0840";
    tmp(40036) := x"0840";
    tmp(40037) := x"001f";
    tmp(40038) := x"001f";
    tmp(40039) := x"001f";
    tmp(40040) := x"001f";
    tmp(40041) := x"001f";
    tmp(40042) := x"001f";
    tmp(40043) := x"001f";
    tmp(40044) := x"001f";
    tmp(40045) := x"001f";
    tmp(40046) := x"001f";
    tmp(40047) := x"001f";
    tmp(40048) := x"001f";
    tmp(40049) := x"001f";
    tmp(40050) := x"001f";
    tmp(40051) := x"001f";
    tmp(40052) := x"001f";
    tmp(40053) := x"001f";
    tmp(40054) := x"001f";
    tmp(40055) := x"001f";
    tmp(40056) := x"001f";
    tmp(40057) := x"001f";
    tmp(40058) := x"001f";
    tmp(40059) := x"001f";
    tmp(40060) := x"001f";
    tmp(40061) := x"001f";
    tmp(40062) := x"001f";
    tmp(40063) := x"001f";
    tmp(40064) := x"001f";
    tmp(40065) := x"001f";
    tmp(40066) := x"001f";
    tmp(40067) := x"001f";
    tmp(40068) := x"001f";
    tmp(40069) := x"001f";
    tmp(40070) := x"001f";
    tmp(40071) := x"001f";
    tmp(40072) := x"001f";
    tmp(40073) := x"001f";
    tmp(40074) := x"001f";
    tmp(40075) := x"001f";
    tmp(40076) := x"001f";
    tmp(40077) := x"1061";
    tmp(40078) := x"1061";
    tmp(40079) := x"1061";
    tmp(40080) := x"0000";
    tmp(40081) := x"0020";
    tmp(40082) := x"0020";
    tmp(40083) := x"0040";
    tmp(40084) := x"0040";
    tmp(40085) := x"0040";
    tmp(40086) := x"0060";
    tmp(40087) := x"0060";
    tmp(40088) := x"0060";
    tmp(40089) := x"0880";
    tmp(40090) := x"0880";
    tmp(40091) := x"08a0";
    tmp(40092) := x"08a0";
    tmp(40093) := x"08a0";
    tmp(40094) := x"08a0";
    tmp(40095) := x"08a0";
    tmp(40096) := x"08a0";
    tmp(40097) := x"08a0";
    tmp(40098) := x"08a0";
    tmp(40099) := x"08c0";
    tmp(40100) := x"08c0";
    tmp(40101) := x"08e0";
    tmp(40102) := x"08e0";
    tmp(40103) := x"08e0";
    tmp(40104) := x"08e0";
    tmp(40105) := x"08e0";
    tmp(40106) := x"0900";
    tmp(40107) := x"0900";
    tmp(40108) := x"0900";
    tmp(40109) := x"0900";
    tmp(40110) := x"0900";
    tmp(40111) := x"0900";
    tmp(40112) := x"0900";
    tmp(40113) := x"0900";
    tmp(40114) := x"1120";
    tmp(40115) := x"1140";
    tmp(40116) := x"1140";
    tmp(40117) := x"1141";
    tmp(40118) := x"1161";
    tmp(40119) := x"1161";
    tmp(40120) := x"1141";
    tmp(40121) := x"1141";
    tmp(40122) := x"1161";
    tmp(40123) := x"1161";
    tmp(40124) := x"1161";
    tmp(40125) := x"1161";
    tmp(40126) := x"1140";
    tmp(40127) := x"1140";
    tmp(40128) := x"1161";
    tmp(40129) := x"1161";
    tmp(40130) := x"1161";
    tmp(40131) := x"1161";
    tmp(40132) := x"1161";
    tmp(40133) := x"1161";
    tmp(40134) := x"1161";
    tmp(40135) := x"1161";
    tmp(40136) := x"1161";
    tmp(40137) := x"1161";
    tmp(40138) := x"1141";
    tmp(40139) := x"1161";
    tmp(40140) := x"1140";
    tmp(40141) := x"1140";
    tmp(40142) := x"1141";
    tmp(40143) := x"1141";
    tmp(40144) := x"1140";
    tmp(40145) := x"1140";
    tmp(40146) := x"1120";
    tmp(40147) := x"0920";
    tmp(40148) := x"0920";
    tmp(40149) := x"0920";
    tmp(40150) := x"0920";
    tmp(40151) := x"0920";
    tmp(40152) := x"0940";
    tmp(40153) := x"1140";
    tmp(40154) := x"0920";
    tmp(40155) := x"0940";
    tmp(40156) := x"0920";
    tmp(40157) := x"0920";
    tmp(40158) := x"0940";
    tmp(40159) := x"0920";
    tmp(40160) := x"0920";
    tmp(40161) := x"0920";
    tmp(40162) := x"0920";
    tmp(40163) := x"0900";
    tmp(40164) := x"0900";
    tmp(40165) := x"0900";
    tmp(40166) := x"0900";
    tmp(40167) := x"0900";
    tmp(40168) := x"0900";
    tmp(40169) := x"0900";
    tmp(40170) := x"0900";
    tmp(40171) := x"0900";
    tmp(40172) := x"0900";
    tmp(40173) := x"0900";
    tmp(40174) := x"0900";
    tmp(40175) := x"0900";
    tmp(40176) := x"0900";
    tmp(40177) := x"0900";
    tmp(40178) := x"0900";
    tmp(40179) := x"0900";
    tmp(40180) := x"0900";
    tmp(40181) := x"0900";
    tmp(40182) := x"0900";
    tmp(40183) := x"0900";
    tmp(40184) := x"0900";
    tmp(40185) := x"0900";
    tmp(40186) := x"0900";
    tmp(40187) := x"08e0";
    tmp(40188) := x"08e0";
    tmp(40189) := x"08e0";
    tmp(40190) := x"08e0";
    tmp(40191) := x"08e0";
    tmp(40192) := x"08e0";
    tmp(40193) := x"08e0";
    tmp(40194) := x"08e0";
    tmp(40195) := x"08c0";
    tmp(40196) := x"08c0";
    tmp(40197) := x"08c0";
    tmp(40198) := x"08c0";
    tmp(40199) := x"08c0";
    tmp(40200) := x"08a0";
    tmp(40201) := x"08a0";
    tmp(40202) := x"08a0";
    tmp(40203) := x"08a0";
    tmp(40204) := x"08a0";
    tmp(40205) := x"08a0";
    tmp(40206) := x"08a0";
    tmp(40207) := x"08a0";
    tmp(40208) := x"08a0";
    tmp(40209) := x"08a0";
    tmp(40210) := x"08a0";
    tmp(40211) := x"08a0";
    tmp(40212) := x"08a0";
    tmp(40213) := x"08c0";
    tmp(40214) := x"08c0";
    tmp(40215) := x"08c0";
    tmp(40216) := x"08c0";
    tmp(40217) := x"08e0";
    tmp(40218) := x"08c0";
    tmp(40219) := x"08c0";
    tmp(40220) := x"08c0";
    tmp(40221) := x"08c0";
    tmp(40222) := x"08c0";
    tmp(40223) := x"08a0";
    tmp(40224) := x"08a0";
    tmp(40225) := x"08a0";
    tmp(40226) := x"08a0";
    tmp(40227) := x"08a0";
    tmp(40228) := x"0880";
    tmp(40229) := x"0880";
    tmp(40230) := x"0860";
    tmp(40231) := x"1060";
    tmp(40232) := x"1060";
    tmp(40233) := x"1060";
    tmp(40234) := x"1060";
    tmp(40235) := x"1060";
    tmp(40236) := x"1060";
    tmp(40237) := x"1060";
    tmp(40238) := x"0860";
    tmp(40239) := x"1840";
    tmp(40240) := x"3840";
    tmp(40241) := x"3040";
    tmp(40242) := x"1840";
    tmp(40243) := x"1840";
    tmp(40244) := x"1840";
    tmp(40245) := x"1840";
    tmp(40246) := x"1840";
    tmp(40247) := x"1040";
    tmp(40248) := x"1040";
    tmp(40249) := x"1040";
    tmp(40250) := x"1040";
    tmp(40251) := x"1040";
    tmp(40252) := x"1040";
    tmp(40253) := x"1040";
    tmp(40254) := x"1040";
    tmp(40255) := x"1040";
    tmp(40256) := x"1060";
    tmp(40257) := x"1040";
    tmp(40258) := x"1061";
    tmp(40259) := x"1060";
    tmp(40260) := x"1060";
    tmp(40261) := x"1061";
    tmp(40262) := x"1061";
    tmp(40263) := x"1061";
    tmp(40264) := x"1061";
    tmp(40265) := x"1061";
    tmp(40266) := x"1060";
    tmp(40267) := x"1060";
    tmp(40268) := x"1040";
    tmp(40269) := x"1040";
    tmp(40270) := x"1040";
    tmp(40271) := x"0840";
    tmp(40272) := x"0840";
    tmp(40273) := x"0840";
    tmp(40274) := x"0840";
    tmp(40275) := x"0840";
    tmp(40276) := x"0840";
    tmp(40277) := x"001f";
    tmp(40278) := x"001f";
    tmp(40279) := x"001f";
    tmp(40280) := x"001f";
    tmp(40281) := x"001f";
    tmp(40282) := x"001f";
    tmp(40283) := x"001f";
    tmp(40284) := x"001f";
    tmp(40285) := x"001f";
    tmp(40286) := x"001f";
    tmp(40287) := x"001f";
    tmp(40288) := x"001f";
    tmp(40289) := x"001f";
    tmp(40290) := x"001f";
    tmp(40291) := x"001f";
    tmp(40292) := x"001f";
    tmp(40293) := x"001f";
    tmp(40294) := x"001f";
    tmp(40295) := x"001f";
    tmp(40296) := x"001f";
    tmp(40297) := x"001f";
    tmp(40298) := x"001f";
    tmp(40299) := x"001f";
    tmp(40300) := x"001f";
    tmp(40301) := x"001f";
    tmp(40302) := x"001f";
    tmp(40303) := x"001f";
    tmp(40304) := x"001f";
    tmp(40305) := x"001f";
    tmp(40306) := x"001f";
    tmp(40307) := x"001f";
    tmp(40308) := x"001f";
    tmp(40309) := x"001f";
    tmp(40310) := x"001f";
    tmp(40311) := x"001f";
    tmp(40312) := x"001f";
    tmp(40313) := x"001f";
    tmp(40314) := x"001f";
    tmp(40315) := x"001f";
    tmp(40316) := x"001f";
    tmp(40317) := x"1061";
    tmp(40318) := x"1061";
    tmp(40319) := x"1061";
    tmp(40320) := x"0000";
    tmp(40321) := x"0040";
    tmp(40322) := x"0040";
    tmp(40323) := x"0040";
    tmp(40324) := x"0060";
    tmp(40325) := x"0060";
    tmp(40326) := x"0060";
    tmp(40327) := x"0060";
    tmp(40328) := x"0060";
    tmp(40329) := x"0880";
    tmp(40330) := x"0880";
    tmp(40331) := x"0880";
    tmp(40332) := x"0880";
    tmp(40333) := x"08a0";
    tmp(40334) := x"08a0";
    tmp(40335) := x"08a0";
    tmp(40336) := x"08a0";
    tmp(40337) := x"08a0";
    tmp(40338) := x"08a0";
    tmp(40339) := x"08a0";
    tmp(40340) := x"08c0";
    tmp(40341) := x"08e0";
    tmp(40342) := x"08e0";
    tmp(40343) := x"08e0";
    tmp(40344) := x"08e0";
    tmp(40345) := x"08e0";
    tmp(40346) := x"08e0";
    tmp(40347) := x"08e0";
    tmp(40348) := x"08e0";
    tmp(40349) := x"0900";
    tmp(40350) := x"0900";
    tmp(40351) := x"0900";
    tmp(40352) := x"0900";
    tmp(40353) := x"0900";
    tmp(40354) := x"0920";
    tmp(40355) := x"1120";
    tmp(40356) := x"1140";
    tmp(40357) := x"1140";
    tmp(40358) := x"1141";
    tmp(40359) := x"1161";
    tmp(40360) := x"1161";
    tmp(40361) := x"1140";
    tmp(40362) := x"1140";
    tmp(40363) := x"1161";
    tmp(40364) := x"1161";
    tmp(40365) := x"1141";
    tmp(40366) := x"1140";
    tmp(40367) := x"1140";
    tmp(40368) := x"1161";
    tmp(40369) := x"1161";
    tmp(40370) := x"1161";
    tmp(40371) := x"1161";
    tmp(40372) := x"1161";
    tmp(40373) := x"1161";
    tmp(40374) := x"1141";
    tmp(40375) := x"1141";
    tmp(40376) := x"1141";
    tmp(40377) := x"1140";
    tmp(40378) := x"1141";
    tmp(40379) := x"1141";
    tmp(40380) := x"1141";
    tmp(40381) := x"1140";
    tmp(40382) := x"1141";
    tmp(40383) := x"1141";
    tmp(40384) := x"1140";
    tmp(40385) := x"1140";
    tmp(40386) := x"0920";
    tmp(40387) := x"0920";
    tmp(40388) := x"0920";
    tmp(40389) := x"0920";
    tmp(40390) := x"0920";
    tmp(40391) := x"0920";
    tmp(40392) := x"0920";
    tmp(40393) := x"0920";
    tmp(40394) := x"0920";
    tmp(40395) := x"0920";
    tmp(40396) := x"0940";
    tmp(40397) := x"0920";
    tmp(40398) := x"0920";
    tmp(40399) := x"0920";
    tmp(40400) := x"0920";
    tmp(40401) := x"0920";
    tmp(40402) := x"0900";
    tmp(40403) := x"0900";
    tmp(40404) := x"0900";
    tmp(40405) := x"0900";
    tmp(40406) := x"0900";
    tmp(40407) := x"0900";
    tmp(40408) := x"0900";
    tmp(40409) := x"0900";
    tmp(40410) := x"0900";
    tmp(40411) := x"0900";
    tmp(40412) := x"0900";
    tmp(40413) := x"0900";
    tmp(40414) := x"0900";
    tmp(40415) := x"0900";
    tmp(40416) := x"0900";
    tmp(40417) := x"0900";
    tmp(40418) := x"0900";
    tmp(40419) := x"0900";
    tmp(40420) := x"0900";
    tmp(40421) := x"0900";
    tmp(40422) := x"0900";
    tmp(40423) := x"0900";
    tmp(40424) := x"0900";
    tmp(40425) := x"08e0";
    tmp(40426) := x"0900";
    tmp(40427) := x"08e0";
    tmp(40428) := x"08e0";
    tmp(40429) := x"08e0";
    tmp(40430) := x"08e0";
    tmp(40431) := x"08e0";
    tmp(40432) := x"08e0";
    tmp(40433) := x"08c0";
    tmp(40434) := x"08c0";
    tmp(40435) := x"08c0";
    tmp(40436) := x"08c0";
    tmp(40437) := x"08c0";
    tmp(40438) := x"08c0";
    tmp(40439) := x"08c0";
    tmp(40440) := x"08a0";
    tmp(40441) := x"08a0";
    tmp(40442) := x"08a0";
    tmp(40443) := x"08a0";
    tmp(40444) := x"08a0";
    tmp(40445) := x"08a0";
    tmp(40446) := x"08a0";
    tmp(40447) := x"08a0";
    tmp(40448) := x"08a0";
    tmp(40449) := x"08a0";
    tmp(40450) := x"08a0";
    tmp(40451) := x"08a0";
    tmp(40452) := x"08a0";
    tmp(40453) := x"08c0";
    tmp(40454) := x"08c0";
    tmp(40455) := x"08c0";
    tmp(40456) := x"08c0";
    tmp(40457) := x"08c0";
    tmp(40458) := x"08c0";
    tmp(40459) := x"08c0";
    tmp(40460) := x"08c0";
    tmp(40461) := x"08c0";
    tmp(40462) := x"08a0";
    tmp(40463) := x"08a0";
    tmp(40464) := x"08a0";
    tmp(40465) := x"08a0";
    tmp(40466) := x"08a0";
    tmp(40467) := x"0880";
    tmp(40468) := x"0880";
    tmp(40469) := x"1080";
    tmp(40470) := x"1060";
    tmp(40471) := x"1060";
    tmp(40472) := x"1060";
    tmp(40473) := x"1060";
    tmp(40474) := x"1060";
    tmp(40475) := x"1060";
    tmp(40476) := x"1040";
    tmp(40477) := x"1040";
    tmp(40478) := x"1040";
    tmp(40479) := x"2020";
    tmp(40480) := x"4020";
    tmp(40481) := x"4020";
    tmp(40482) := x"3820";
    tmp(40483) := x"3020";
    tmp(40484) := x"4840";
    tmp(40485) := x"5040";
    tmp(40486) := x"5041";
    tmp(40487) := x"3841";
    tmp(40488) := x"2061";
    tmp(40489) := x"1040";
    tmp(40490) := x"1040";
    tmp(40491) := x"1040";
    tmp(40492) := x"1040";
    tmp(40493) := x"1040";
    tmp(40494) := x"1040";
    tmp(40495) := x"1040";
    tmp(40496) := x"1040";
    tmp(40497) := x"1040";
    tmp(40498) := x"1060";
    tmp(40499) := x"1060";
    tmp(40500) := x"1060";
    tmp(40501) := x"1060";
    tmp(40502) := x"1060";
    tmp(40503) := x"1061";
    tmp(40504) := x"1061";
    tmp(40505) := x"1060";
    tmp(40506) := x"1060";
    tmp(40507) := x"1060";
    tmp(40508) := x"1040";
    tmp(40509) := x"1040";
    tmp(40510) := x"0840";
    tmp(40511) := x"0840";
    tmp(40512) := x"0840";
    tmp(40513) := x"0840";
    tmp(40514) := x"0840";
    tmp(40515) := x"0840";
    tmp(40516) := x"0840";
    tmp(40517) := x"001f";
    tmp(40518) := x"001f";
    tmp(40519) := x"001f";
    tmp(40520) := x"001f";
    tmp(40521) := x"001f";
    tmp(40522) := x"001f";
    tmp(40523) := x"001f";
    tmp(40524) := x"001f";
    tmp(40525) := x"001f";
    tmp(40526) := x"001f";
    tmp(40527) := x"001f";
    tmp(40528) := x"001f";
    tmp(40529) := x"001f";
    tmp(40530) := x"001f";
    tmp(40531) := x"001f";
    tmp(40532) := x"001f";
    tmp(40533) := x"001f";
    tmp(40534) := x"001f";
    tmp(40535) := x"001f";
    tmp(40536) := x"001f";
    tmp(40537) := x"001f";
    tmp(40538) := x"001f";
    tmp(40539) := x"001f";
    tmp(40540) := x"001f";
    tmp(40541) := x"001f";
    tmp(40542) := x"001f";
    tmp(40543) := x"001f";
    tmp(40544) := x"001f";
    tmp(40545) := x"001f";
    tmp(40546) := x"001f";
    tmp(40547) := x"001f";
    tmp(40548) := x"001f";
    tmp(40549) := x"001f";
    tmp(40550) := x"001f";
    tmp(40551) := x"001f";
    tmp(40552) := x"001f";
    tmp(40553) := x"001f";
    tmp(40554) := x"001f";
    tmp(40555) := x"001f";
    tmp(40556) := x"001f";
    tmp(40557) := x"1061";
    tmp(40558) := x"1061";
    tmp(40559) := x"1061";
    tmp(40560) := x"0000";
    tmp(40561) := x"0060";
    tmp(40562) := x"0040";
    tmp(40563) := x"0040";
    tmp(40564) := x"0060";
    tmp(40565) := x"0060";
    tmp(40566) := x"0060";
    tmp(40567) := x"0060";
    tmp(40568) := x"0860";
    tmp(40569) := x"0860";
    tmp(40570) := x"0860";
    tmp(40571) := x"0880";
    tmp(40572) := x"0880";
    tmp(40573) := x"0880";
    tmp(40574) := x"0880";
    tmp(40575) := x"0880";
    tmp(40576) := x"08a0";
    tmp(40577) := x"08a0";
    tmp(40578) := x"08a0";
    tmp(40579) := x"08a0";
    tmp(40580) := x"08a0";
    tmp(40581) := x"08c0";
    tmp(40582) := x"08c0";
    tmp(40583) := x"08e0";
    tmp(40584) := x"08e0";
    tmp(40585) := x"08e0";
    tmp(40586) := x"08e0";
    tmp(40587) := x"08e0";
    tmp(40588) := x"08e0";
    tmp(40589) := x"08e0";
    tmp(40590) := x"0900";
    tmp(40591) := x"0900";
    tmp(40592) := x"0900";
    tmp(40593) := x"0900";
    tmp(40594) := x"0900";
    tmp(40595) := x"0920";
    tmp(40596) := x"1120";
    tmp(40597) := x"1140";
    tmp(40598) := x"1141";
    tmp(40599) := x"1141";
    tmp(40600) := x"1140";
    tmp(40601) := x"1141";
    tmp(40602) := x"1140";
    tmp(40603) := x"1140";
    tmp(40604) := x"1140";
    tmp(40605) := x"1141";
    tmp(40606) := x"1140";
    tmp(40607) := x"1140";
    tmp(40608) := x"1161";
    tmp(40609) := x"1161";
    tmp(40610) := x"1181";
    tmp(40611) := x"1181";
    tmp(40612) := x"1161";
    tmp(40613) := x"1161";
    tmp(40614) := x"1141";
    tmp(40615) := x"1141";
    tmp(40616) := x"1141";
    tmp(40617) := x"1141";
    tmp(40618) := x"1141";
    tmp(40619) := x"1141";
    tmp(40620) := x"1141";
    tmp(40621) := x"1140";
    tmp(40622) := x"1141";
    tmp(40623) := x"1141";
    tmp(40624) := x"1140";
    tmp(40625) := x"1140";
    tmp(40626) := x"0920";
    tmp(40627) := x"0920";
    tmp(40628) := x"0920";
    tmp(40629) := x"0920";
    tmp(40630) := x"0920";
    tmp(40631) := x"0920";
    tmp(40632) := x"0920";
    tmp(40633) := x"0920";
    tmp(40634) := x"0920";
    tmp(40635) := x"0920";
    tmp(40636) := x"0920";
    tmp(40637) := x"0920";
    tmp(40638) := x"0920";
    tmp(40639) := x"0920";
    tmp(40640) := x"0920";
    tmp(40641) := x"0920";
    tmp(40642) := x"0920";
    tmp(40643) := x"0900";
    tmp(40644) := x"0900";
    tmp(40645) := x"0900";
    tmp(40646) := x"0900";
    tmp(40647) := x"0900";
    tmp(40648) := x"0900";
    tmp(40649) := x"0900";
    tmp(40650) := x"0900";
    tmp(40651) := x"0900";
    tmp(40652) := x"0900";
    tmp(40653) := x"0900";
    tmp(40654) := x"0900";
    tmp(40655) := x"0900";
    tmp(40656) := x"0900";
    tmp(40657) := x"0900";
    tmp(40658) := x"0900";
    tmp(40659) := x"0900";
    tmp(40660) := x"0900";
    tmp(40661) := x"0900";
    tmp(40662) := x"0900";
    tmp(40663) := x"0900";
    tmp(40664) := x"08e0";
    tmp(40665) := x"0900";
    tmp(40666) := x"0900";
    tmp(40667) := x"0900";
    tmp(40668) := x"08e0";
    tmp(40669) := x"08e0";
    tmp(40670) := x"08e0";
    tmp(40671) := x"08e0";
    tmp(40672) := x"08c0";
    tmp(40673) := x"08c0";
    tmp(40674) := x"08c0";
    tmp(40675) := x"08c0";
    tmp(40676) := x"08c0";
    tmp(40677) := x"08c0";
    tmp(40678) := x"08c0";
    tmp(40679) := x"08a0";
    tmp(40680) := x"08a0";
    tmp(40681) := x"08a0";
    tmp(40682) := x"08a0";
    tmp(40683) := x"08a0";
    tmp(40684) := x"08a0";
    tmp(40685) := x"08a0";
    tmp(40686) := x"08a0";
    tmp(40687) := x"08a0";
    tmp(40688) := x"08a0";
    tmp(40689) := x"08a0";
    tmp(40690) := x"08a0";
    tmp(40691) := x"08a0";
    tmp(40692) := x"0880";
    tmp(40693) := x"0880";
    tmp(40694) := x"0880";
    tmp(40695) := x"0880";
    tmp(40696) := x"0880";
    tmp(40697) := x"0880";
    tmp(40698) := x"0880";
    tmp(40699) := x"0880";
    tmp(40700) := x"0880";
    tmp(40701) := x"0880";
    tmp(40702) := x"0880";
    tmp(40703) := x"0880";
    tmp(40704) := x"0860";
    tmp(40705) := x"0860";
    tmp(40706) := x"0860";
    tmp(40707) := x"0860";
    tmp(40708) := x"0880";
    tmp(40709) := x"1080";
    tmp(40710) := x"1060";
    tmp(40711) := x"1060";
    tmp(40712) := x"1060";
    tmp(40713) := x"1060";
    tmp(40714) := x"1060";
    tmp(40715) := x"1060";
    tmp(40716) := x"1040";
    tmp(40717) := x"1840";
    tmp(40718) := x"2020";
    tmp(40719) := x"2800";
    tmp(40720) := x"3000";
    tmp(40721) := x"3000";
    tmp(40722) := x"4000";
    tmp(40723) := x"4800";
    tmp(40724) := x"6820";
    tmp(40725) := x"6820";
    tmp(40726) := x"7820";
    tmp(40727) := x"8020";
    tmp(40728) := x"6841";
    tmp(40729) := x"3841";
    tmp(40730) := x"1840";
    tmp(40731) := x"1040";
    tmp(40732) := x"1040";
    tmp(40733) := x"1060";
    tmp(40734) := x"1060";
    tmp(40735) := x"1060";
    tmp(40736) := x"1060";
    tmp(40737) := x"1060";
    tmp(40738) := x"1060";
    tmp(40739) := x"1060";
    tmp(40740) := x"1060";
    tmp(40741) := x"1060";
    tmp(40742) := x"1061";
    tmp(40743) := x"1061";
    tmp(40744) := x"1061";
    tmp(40745) := x"1060";
    tmp(40746) := x"1060";
    tmp(40747) := x"1060";
    tmp(40748) := x"1040";
    tmp(40749) := x"1040";
    tmp(40750) := x"0840";
    tmp(40751) := x"0840";
    tmp(40752) := x"0840";
    tmp(40753) := x"0840";
    tmp(40754) := x"0840";
    tmp(40755) := x"0840";
    tmp(40756) := x"0840";
    tmp(40757) := x"001f";
    tmp(40758) := x"001f";
    tmp(40759) := x"001f";
    tmp(40760) := x"001f";
    tmp(40761) := x"001f";
    tmp(40762) := x"001f";
    tmp(40763) := x"001f";
    tmp(40764) := x"001f";
    tmp(40765) := x"001f";
    tmp(40766) := x"001f";
    tmp(40767) := x"001f";
    tmp(40768) := x"001f";
    tmp(40769) := x"001f";
    tmp(40770) := x"001f";
    tmp(40771) := x"001f";
    tmp(40772) := x"001f";
    tmp(40773) := x"001f";
    tmp(40774) := x"001f";
    tmp(40775) := x"001f";
    tmp(40776) := x"001f";
    tmp(40777) := x"001f";
    tmp(40778) := x"001f";
    tmp(40779) := x"001f";
    tmp(40780) := x"001f";
    tmp(40781) := x"001f";
    tmp(40782) := x"001f";
    tmp(40783) := x"001f";
    tmp(40784) := x"001f";
    tmp(40785) := x"001f";
    tmp(40786) := x"001f";
    tmp(40787) := x"001f";
    tmp(40788) := x"001f";
    tmp(40789) := x"001f";
    tmp(40790) := x"001f";
    tmp(40791) := x"001f";
    tmp(40792) := x"001f";
    tmp(40793) := x"001f";
    tmp(40794) := x"001f";
    tmp(40795) := x"001f";
    tmp(40796) := x"001f";
    tmp(40797) := x"1061";
    tmp(40798) := x"1061";
    tmp(40799) := x"1061";
    tmp(40800) := x"0000";
    tmp(40801) := x"0040";
    tmp(40802) := x"0040";
    tmp(40803) := x"0040";
    tmp(40804) := x"0860";
    tmp(40805) := x"0040";
    tmp(40806) := x"0860";
    tmp(40807) := x"0060";
    tmp(40808) := x"0860";
    tmp(40809) := x"0860";
    tmp(40810) := x"0860";
    tmp(40811) := x"0860";
    tmp(40812) := x"0880";
    tmp(40813) := x"0880";
    tmp(40814) := x"0880";
    tmp(40815) := x"0880";
    tmp(40816) := x"0880";
    tmp(40817) := x"0880";
    tmp(40818) := x"08a0";
    tmp(40819) := x"08a0";
    tmp(40820) := x"08a0";
    tmp(40821) := x"08a0";
    tmp(40822) := x"08c0";
    tmp(40823) := x"08c0";
    tmp(40824) := x"08c0";
    tmp(40825) := x"08c0";
    tmp(40826) := x"08c0";
    tmp(40827) := x"08e0";
    tmp(40828) := x"08e0";
    tmp(40829) := x"08e0";
    tmp(40830) := x"08e0";
    tmp(40831) := x"0900";
    tmp(40832) := x"0900";
    tmp(40833) := x"0900";
    tmp(40834) := x"0900";
    tmp(40835) := x"0920";
    tmp(40836) := x"1120";
    tmp(40837) := x"1120";
    tmp(40838) := x"1140";
    tmp(40839) := x"1140";
    tmp(40840) := x"1140";
    tmp(40841) := x"1140";
    tmp(40842) := x"1140";
    tmp(40843) := x"1120";
    tmp(40844) := x"1140";
    tmp(40845) := x"1140";
    tmp(40846) := x"1140";
    tmp(40847) := x"1140";
    tmp(40848) := x"1141";
    tmp(40849) := x"1161";
    tmp(40850) := x"1161";
    tmp(40851) := x"1181";
    tmp(40852) := x"1161";
    tmp(40853) := x"1161";
    tmp(40854) := x"1141";
    tmp(40855) := x"1141";
    tmp(40856) := x"1141";
    tmp(40857) := x"1141";
    tmp(40858) := x"1141";
    tmp(40859) := x"1141";
    tmp(40860) := x"1141";
    tmp(40861) := x"1141";
    tmp(40862) := x"1140";
    tmp(40863) := x"1140";
    tmp(40864) := x"1140";
    tmp(40865) := x"1120";
    tmp(40866) := x"0920";
    tmp(40867) := x"0920";
    tmp(40868) := x"0920";
    tmp(40869) := x"0920";
    tmp(40870) := x"0920";
    tmp(40871) := x"0920";
    tmp(40872) := x"0920";
    tmp(40873) := x"0920";
    tmp(40874) := x"0920";
    tmp(40875) := x"0920";
    tmp(40876) := x"0920";
    tmp(40877) := x"0920";
    tmp(40878) := x"0920";
    tmp(40879) := x"0920";
    tmp(40880) := x"0920";
    tmp(40881) := x"0920";
    tmp(40882) := x"0900";
    tmp(40883) := x"0900";
    tmp(40884) := x"0900";
    tmp(40885) := x"0900";
    tmp(40886) := x"0900";
    tmp(40887) := x"08e0";
    tmp(40888) := x"0900";
    tmp(40889) := x"0900";
    tmp(40890) := x"0900";
    tmp(40891) := x"0900";
    tmp(40892) := x"0900";
    tmp(40893) := x"0900";
    tmp(40894) := x"0900";
    tmp(40895) := x"0900";
    tmp(40896) := x"0900";
    tmp(40897) := x"0900";
    tmp(40898) := x"0900";
    tmp(40899) := x"0900";
    tmp(40900) := x"0900";
    tmp(40901) := x"0900";
    tmp(40902) := x"0900";
    tmp(40903) := x"0900";
    tmp(40904) := x"0900";
    tmp(40905) := x"0900";
    tmp(40906) := x"08e0";
    tmp(40907) := x"08e0";
    tmp(40908) := x"08e0";
    tmp(40909) := x"08e0";
    tmp(40910) := x"08e0";
    tmp(40911) := x"08e0";
    tmp(40912) := x"08c0";
    tmp(40913) := x"08c0";
    tmp(40914) := x"08c0";
    tmp(40915) := x"08c0";
    tmp(40916) := x"08c0";
    tmp(40917) := x"08a0";
    tmp(40918) := x"08c0";
    tmp(40919) := x"08a0";
    tmp(40920) := x"08a0";
    tmp(40921) := x"08a0";
    tmp(40922) := x"08a0";
    tmp(40923) := x"08a0";
    tmp(40924) := x"08a0";
    tmp(40925) := x"08a0";
    tmp(40926) := x"08a0";
    tmp(40927) := x"0880";
    tmp(40928) := x"0860";
    tmp(40929) := x"0860";
    tmp(40930) := x"0880";
    tmp(40931) := x"10a0";
    tmp(40932) := x"1901";
    tmp(40933) := x"2981";
    tmp(40934) := x"4222";
    tmp(40935) := x"4a42";
    tmp(40936) := x"5263";
    tmp(40937) := x"5a83";
    tmp(40938) := x"62a3";
    tmp(40939) := x"5a83";
    tmp(40940) := x"6283";
    tmp(40941) := x"7b65";
    tmp(40942) := x"8be7";
    tmp(40943) := x"8366";
    tmp(40944) := x"7345";
    tmp(40945) := x"5aa4";
    tmp(40946) := x"4203";
    tmp(40947) := x"2921";
    tmp(40948) := x"18a1";
    tmp(40949) := x"0860";
    tmp(40950) := x"0840";
    tmp(40951) := x"0840";
    tmp(40952) := x"1060";
    tmp(40953) := x"1060";
    tmp(40954) := x"1060";
    tmp(40955) := x"1060";
    tmp(40956) := x"1840";
    tmp(40957) := x"2820";
    tmp(40958) := x"2000";
    tmp(40959) := x"2800";
    tmp(40960) := x"2800";
    tmp(40961) := x"2800";
    tmp(40962) := x"3800";
    tmp(40963) := x"5000";
    tmp(40964) := x"5800";
    tmp(40965) := x"5000";
    tmp(40966) := x"6800";
    tmp(40967) := x"9020";
    tmp(40968) := x"9020";
    tmp(40969) := x"6841";
    tmp(40970) := x"3061";
    tmp(40971) := x"1040";
    tmp(40972) := x"1040";
    tmp(40973) := x"1040";
    tmp(40974) := x"1040";
    tmp(40975) := x"1040";
    tmp(40976) := x"1040";
    tmp(40977) := x"1040";
    tmp(40978) := x"1060";
    tmp(40979) := x"1060";
    tmp(40980) := x"1060";
    tmp(40981) := x"1060";
    tmp(40982) := x"1061";
    tmp(40983) := x"1061";
    tmp(40984) := x"1060";
    tmp(40985) := x"1060";
    tmp(40986) := x"1060";
    tmp(40987) := x"1040";
    tmp(40988) := x"1040";
    tmp(40989) := x"0840";
    tmp(40990) := x"0840";
    tmp(40991) := x"0840";
    tmp(40992) := x"0840";
    tmp(40993) := x"0840";
    tmp(40994) := x"0840";
    tmp(40995) := x"0840";
    tmp(40996) := x"0840";
    tmp(40997) := x"001f";
    tmp(40998) := x"001f";
    tmp(40999) := x"001f";
    tmp(41000) := x"001f";
    tmp(41001) := x"001f";
    tmp(41002) := x"001f";
    tmp(41003) := x"001f";
    tmp(41004) := x"001f";
    tmp(41005) := x"001f";
    tmp(41006) := x"001f";
    tmp(41007) := x"001f";
    tmp(41008) := x"001f";
    tmp(41009) := x"001f";
    tmp(41010) := x"001f";
    tmp(41011) := x"001f";
    tmp(41012) := x"001f";
    tmp(41013) := x"001f";
    tmp(41014) := x"001f";
    tmp(41015) := x"001f";
    tmp(41016) := x"001f";
    tmp(41017) := x"001f";
    tmp(41018) := x"001f";
    tmp(41019) := x"001f";
    tmp(41020) := x"001f";
    tmp(41021) := x"001f";
    tmp(41022) := x"001f";
    tmp(41023) := x"001f";
    tmp(41024) := x"001f";
    tmp(41025) := x"001f";
    tmp(41026) := x"001f";
    tmp(41027) := x"001f";
    tmp(41028) := x"001f";
    tmp(41029) := x"001f";
    tmp(41030) := x"001f";
    tmp(41031) := x"001f";
    tmp(41032) := x"001f";
    tmp(41033) := x"001f";
    tmp(41034) := x"001f";
    tmp(41035) := x"001f";
    tmp(41036) := x"001f";
    tmp(41037) := x"1061";
    tmp(41038) := x"1061";
    tmp(41039) := x"1061";
    tmp(41040) := x"0000";
    tmp(41041) := x"0860";
    tmp(41042) := x"0860";
    tmp(41043) := x"0840";
    tmp(41044) := x"0840";
    tmp(41045) := x"0840";
    tmp(41046) := x"0840";
    tmp(41047) := x"0860";
    tmp(41048) := x"0860";
    tmp(41049) := x"0860";
    tmp(41050) := x"0860";
    tmp(41051) := x"0860";
    tmp(41052) := x"0860";
    tmp(41053) := x"0860";
    tmp(41054) := x"0880";
    tmp(41055) := x"0880";
    tmp(41056) := x"0880";
    tmp(41057) := x"0880";
    tmp(41058) := x"0880";
    tmp(41059) := x"08a0";
    tmp(41060) := x"08a0";
    tmp(41061) := x"08a0";
    tmp(41062) := x"08a0";
    tmp(41063) := x"08c0";
    tmp(41064) := x"08c0";
    tmp(41065) := x"08c0";
    tmp(41066) := x"08c0";
    tmp(41067) := x"08c0";
    tmp(41068) := x"08e0";
    tmp(41069) := x"08e0";
    tmp(41070) := x"08e0";
    tmp(41071) := x"0900";
    tmp(41072) := x"08e0";
    tmp(41073) := x"0900";
    tmp(41074) := x"0900";
    tmp(41075) := x"0900";
    tmp(41076) := x"0920";
    tmp(41077) := x"0920";
    tmp(41078) := x"1120";
    tmp(41079) := x"1140";
    tmp(41080) := x"1140";
    tmp(41081) := x"1140";
    tmp(41082) := x"1140";
    tmp(41083) := x"1140";
    tmp(41084) := x"1140";
    tmp(41085) := x"1120";
    tmp(41086) := x"1140";
    tmp(41087) := x"1140";
    tmp(41088) := x"1140";
    tmp(41089) := x"1160";
    tmp(41090) := x"1161";
    tmp(41091) := x"1161";
    tmp(41092) := x"1181";
    tmp(41093) := x"1161";
    tmp(41094) := x"1161";
    tmp(41095) := x"1161";
    tmp(41096) := x"1141";
    tmp(41097) := x"1141";
    tmp(41098) := x"1140";
    tmp(41099) := x"1141";
    tmp(41100) := x"1120";
    tmp(41101) := x"1120";
    tmp(41102) := x"1141";
    tmp(41103) := x"1140";
    tmp(41104) := x"1140";
    tmp(41105) := x"1140";
    tmp(41106) := x"0920";
    tmp(41107) := x"0920";
    tmp(41108) := x"0920";
    tmp(41109) := x"0920";
    tmp(41110) := x"0900";
    tmp(41111) := x"0920";
    tmp(41112) := x"0920";
    tmp(41113) := x"0920";
    tmp(41114) := x"0940";
    tmp(41115) := x"0940";
    tmp(41116) := x"0920";
    tmp(41117) := x"0920";
    tmp(41118) := x"0920";
    tmp(41119) := x"0920";
    tmp(41120) := x"0920";
    tmp(41121) := x"0920";
    tmp(41122) := x"0900";
    tmp(41123) := x"0900";
    tmp(41124) := x"0900";
    tmp(41125) := x"0900";
    tmp(41126) := x"0900";
    tmp(41127) := x"08e0";
    tmp(41128) := x"0900";
    tmp(41129) := x"0900";
    tmp(41130) := x"0900";
    tmp(41131) := x"0900";
    tmp(41132) := x"0900";
    tmp(41133) := x"0900";
    tmp(41134) := x"0900";
    tmp(41135) := x"0900";
    tmp(41136) := x"0900";
    tmp(41137) := x"0900";
    tmp(41138) := x"0920";
    tmp(41139) := x"0920";
    tmp(41140) := x"0900";
    tmp(41141) := x"0900";
    tmp(41142) := x"0900";
    tmp(41143) := x"0900";
    tmp(41144) := x"0900";
    tmp(41145) := x"0900";
    tmp(41146) := x"08e0";
    tmp(41147) := x"08e0";
    tmp(41148) := x"08e0";
    tmp(41149) := x"08e0";
    tmp(41150) := x"08e0";
    tmp(41151) := x"08c0";
    tmp(41152) := x"08c0";
    tmp(41153) := x"08c0";
    tmp(41154) := x"08c0";
    tmp(41155) := x"08c0";
    tmp(41156) := x"08c0";
    tmp(41157) := x"08a0";
    tmp(41158) := x"08a0";
    tmp(41159) := x"08a0";
    tmp(41160) := x"08a0";
    tmp(41161) := x"08a0";
    tmp(41162) := x"08a0";
    tmp(41163) := x"08a0";
    tmp(41164) := x"08a0";
    tmp(41165) := x"0880";
    tmp(41166) := x"0880";
    tmp(41167) := x"18e0";
    tmp(41168) := x"31a2";
    tmp(41169) := x"62a4";
    tmp(41170) := x"7b26";
    tmp(41171) := x"9387";
    tmp(41172) := x"ac09";
    tmp(41173) := x"b40a";
    tmp(41174) := x"cc8b";
    tmp(41175) := x"d4ec";
    tmp(41176) := x"e4ec";
    tmp(41177) := x"d44b";
    tmp(41178) := x"c3c9";
    tmp(41179) := x"cbea";
    tmp(41180) := x"ed2d";
    tmp(41181) := x"fdae";
    tmp(41182) := x"ed2d";
    tmp(41183) := x"ed0d";
    tmp(41184) := x"fd6e";
    tmp(41185) := x"f58e";
    tmp(41186) := x"e56d";
    tmp(41187) := x"d54d";
    tmp(41188) := x"bd6d";
    tmp(41189) := x"a46b";
    tmp(41190) := x"6ac7";
    tmp(41191) := x"4163";
    tmp(41192) := x"1881";
    tmp(41193) := x"0840";
    tmp(41194) := x"0840";
    tmp(41195) := x"1040";
    tmp(41196) := x"2040";
    tmp(41197) := x"2000";
    tmp(41198) := x"1800";
    tmp(41199) := x"2000";
    tmp(41200) := x"2000";
    tmp(41201) := x"2800";
    tmp(41202) := x"3000";
    tmp(41203) := x"4000";
    tmp(41204) := x"4000";
    tmp(41205) := x"4800";
    tmp(41206) := x"5800";
    tmp(41207) := x"6800";
    tmp(41208) := x"7020";
    tmp(41209) := x"8020";
    tmp(41210) := x"7041";
    tmp(41211) := x"4061";
    tmp(41212) := x"1840";
    tmp(41213) := x"1040";
    tmp(41214) := x"1040";
    tmp(41215) := x"1040";
    tmp(41216) := x"1040";
    tmp(41217) := x"1040";
    tmp(41218) := x"1040";
    tmp(41219) := x"1040";
    tmp(41220) := x"1040";
    tmp(41221) := x"1060";
    tmp(41222) := x"1060";
    tmp(41223) := x"1060";
    tmp(41224) := x"1040";
    tmp(41225) := x"1040";
    tmp(41226) := x"1060";
    tmp(41227) := x"1040";
    tmp(41228) := x"1040";
    tmp(41229) := x"0840";
    tmp(41230) := x"0840";
    tmp(41231) := x"0840";
    tmp(41232) := x"0840";
    tmp(41233) := x"0840";
    tmp(41234) := x"0840";
    tmp(41235) := x"0840";
    tmp(41236) := x"0840";
    tmp(41237) := x"001f";
    tmp(41238) := x"001f";
    tmp(41239) := x"001f";
    tmp(41240) := x"001f";
    tmp(41241) := x"001f";
    tmp(41242) := x"001f";
    tmp(41243) := x"001f";
    tmp(41244) := x"001f";
    tmp(41245) := x"001f";
    tmp(41246) := x"001f";
    tmp(41247) := x"001f";
    tmp(41248) := x"001f";
    tmp(41249) := x"001f";
    tmp(41250) := x"001f";
    tmp(41251) := x"001f";
    tmp(41252) := x"001f";
    tmp(41253) := x"001f";
    tmp(41254) := x"001f";
    tmp(41255) := x"001f";
    tmp(41256) := x"001f";
    tmp(41257) := x"001f";
    tmp(41258) := x"001f";
    tmp(41259) := x"001f";
    tmp(41260) := x"001f";
    tmp(41261) := x"001f";
    tmp(41262) := x"001f";
    tmp(41263) := x"001f";
    tmp(41264) := x"001f";
    tmp(41265) := x"001f";
    tmp(41266) := x"001f";
    tmp(41267) := x"001f";
    tmp(41268) := x"001f";
    tmp(41269) := x"001f";
    tmp(41270) := x"001f";
    tmp(41271) := x"001f";
    tmp(41272) := x"001f";
    tmp(41273) := x"001f";
    tmp(41274) := x"001f";
    tmp(41275) := x"001f";
    tmp(41276) := x"001f";
    tmp(41277) := x"1061";
    tmp(41278) := x"1061";
    tmp(41279) := x"1061";
    tmp(41280) := x"0000";
    tmp(41281) := x"0860";
    tmp(41282) := x"0860";
    tmp(41283) := x"0840";
    tmp(41284) := x"0860";
    tmp(41285) := x"0840";
    tmp(41286) := x"0840";
    tmp(41287) := x"0860";
    tmp(41288) := x"0860";
    tmp(41289) := x"0860";
    tmp(41290) := x"0860";
    tmp(41291) := x"0860";
    tmp(41292) := x"0860";
    tmp(41293) := x"0860";
    tmp(41294) := x"0860";
    tmp(41295) := x"0880";
    tmp(41296) := x"0880";
    tmp(41297) := x"0880";
    tmp(41298) := x"0880";
    tmp(41299) := x"0880";
    tmp(41300) := x"0880";
    tmp(41301) := x"0880";
    tmp(41302) := x"08a0";
    tmp(41303) := x"08a0";
    tmp(41304) := x"08a0";
    tmp(41305) := x"08c0";
    tmp(41306) := x"08c0";
    tmp(41307) := x"08c0";
    tmp(41308) := x"08c0";
    tmp(41309) := x"08c0";
    tmp(41310) := x"08e0";
    tmp(41311) := x"08e0";
    tmp(41312) := x"0900";
    tmp(41313) := x"0900";
    tmp(41314) := x"0900";
    tmp(41315) := x"0900";
    tmp(41316) := x"0900";
    tmp(41317) := x"0920";
    tmp(41318) := x"0920";
    tmp(41319) := x"1120";
    tmp(41320) := x"1140";
    tmp(41321) := x"1140";
    tmp(41322) := x"1140";
    tmp(41323) := x"1140";
    tmp(41324) := x"1120";
    tmp(41325) := x"1140";
    tmp(41326) := x"1140";
    tmp(41327) := x"1140";
    tmp(41328) := x"1140";
    tmp(41329) := x"1140";
    tmp(41330) := x"1160";
    tmp(41331) := x"1161";
    tmp(41332) := x"1161";
    tmp(41333) := x"1161";
    tmp(41334) := x"1161";
    tmp(41335) := x"1141";
    tmp(41336) := x"1141";
    tmp(41337) := x"1141";
    tmp(41338) := x"1140";
    tmp(41339) := x"1141";
    tmp(41340) := x"1141";
    tmp(41341) := x"1141";
    tmp(41342) := x"1141";
    tmp(41343) := x"1140";
    tmp(41344) := x"1140";
    tmp(41345) := x"1120";
    tmp(41346) := x"0920";
    tmp(41347) := x"0920";
    tmp(41348) := x"0920";
    tmp(41349) := x"0920";
    tmp(41350) := x"0920";
    tmp(41351) := x"0920";
    tmp(41352) := x"0920";
    tmp(41353) := x"0920";
    tmp(41354) := x"0940";
    tmp(41355) := x"0920";
    tmp(41356) := x"0940";
    tmp(41357) := x"0920";
    tmp(41358) := x"0920";
    tmp(41359) := x"0920";
    tmp(41360) := x"0920";
    tmp(41361) := x"0920";
    tmp(41362) := x"0920";
    tmp(41363) := x"0900";
    tmp(41364) := x"0900";
    tmp(41365) := x"0900";
    tmp(41366) := x"0900";
    tmp(41367) := x"0900";
    tmp(41368) := x"0900";
    tmp(41369) := x"0900";
    tmp(41370) := x"0900";
    tmp(41371) := x"0900";
    tmp(41372) := x"0900";
    tmp(41373) := x"0900";
    tmp(41374) := x"0900";
    tmp(41375) := x"0900";
    tmp(41376) := x"0920";
    tmp(41377) := x"0900";
    tmp(41378) := x"0920";
    tmp(41379) := x"0920";
    tmp(41380) := x"0900";
    tmp(41381) := x"0900";
    tmp(41382) := x"0900";
    tmp(41383) := x"0900";
    tmp(41384) := x"0900";
    tmp(41385) := x"0900";
    tmp(41386) := x"0900";
    tmp(41387) := x"08e0";
    tmp(41388) := x"0900";
    tmp(41389) := x"08e0";
    tmp(41390) := x"08e0";
    tmp(41391) := x"08c0";
    tmp(41392) := x"08c0";
    tmp(41393) := x"08c0";
    tmp(41394) := x"08c0";
    tmp(41395) := x"08c0";
    tmp(41396) := x"08c0";
    tmp(41397) := x"08c0";
    tmp(41398) := x"08a0";
    tmp(41399) := x"08a0";
    tmp(41400) := x"08a0";
    tmp(41401) := x"08a0";
    tmp(41402) := x"0880";
    tmp(41403) := x"0860";
    tmp(41404) := x"10c0";
    tmp(41405) := x"41e2";
    tmp(41406) := x"8b66";
    tmp(41407) := x"b3e9";
    tmp(41408) := x"bbea";
    tmp(41409) := x"c3eb";
    tmp(41410) := x"d46c";
    tmp(41411) := x"dc8d";
    tmp(41412) := x"d44d";
    tmp(41413) := x"dc6d";
    tmp(41414) := x"ecce";
    tmp(41415) := x"fdb0";
    tmp(41416) := x"fdb1";
    tmp(41417) := x"ecce";
    tmp(41418) := x"cbaa";
    tmp(41419) := x"e42b";
    tmp(41420) := x"f4ee";
    tmp(41421) := x"fd6f";
    tmp(41422) := x"f52e";
    tmp(41423) := x"f4ee";
    tmp(41424) := x"f4ee";
    tmp(41425) := x"fd4f";
    tmp(41426) := x"fdb1";
    tmp(41427) := x"fd50";
    tmp(41428) := x"fe13";
    tmp(41429) := x"fdf3";
    tmp(41430) := x"f5f3";
    tmp(41431) := x"e653";
    tmp(41432) := x"d634";
    tmp(41433) := x"a44d";
    tmp(41434) := x"49e5";
    tmp(41435) := x"2081";
    tmp(41436) := x"2040";
    tmp(41437) := x"2000";
    tmp(41438) := x"1800";
    tmp(41439) := x"1800";
    tmp(41440) := x"1800";
    tmp(41441) := x"2000";
    tmp(41442) := x"3000";
    tmp(41443) := x"3800";
    tmp(41444) := x"3800";
    tmp(41445) := x"3000";
    tmp(41446) := x"4800";
    tmp(41447) := x"5000";
    tmp(41448) := x"5000";
    tmp(41449) := x"8020";
    tmp(41450) := x"a841";
    tmp(41451) := x"b061";
    tmp(41452) := x"5061";
    tmp(41453) := x"1840";
    tmp(41454) := x"1040";
    tmp(41455) := x"1040";
    tmp(41456) := x"1060";
    tmp(41457) := x"1040";
    tmp(41458) := x"1040";
    tmp(41459) := x"1061";
    tmp(41460) := x"1040";
    tmp(41461) := x"1040";
    tmp(41462) := x"1060";
    tmp(41463) := x"1060";
    tmp(41464) := x"1060";
    tmp(41465) := x"1060";
    tmp(41466) := x"1040";
    tmp(41467) := x"1040";
    tmp(41468) := x"0840";
    tmp(41469) := x"0840";
    tmp(41470) := x"0840";
    tmp(41471) := x"0840";
    tmp(41472) := x"0840";
    tmp(41473) := x"0840";
    tmp(41474) := x"0840";
    tmp(41475) := x"0840";
    tmp(41476) := x"0840";
    tmp(41477) := x"001f";
    tmp(41478) := x"001f";
    tmp(41479) := x"001f";
    tmp(41480) := x"001f";
    tmp(41481) := x"001f";
    tmp(41482) := x"001f";
    tmp(41483) := x"001f";
    tmp(41484) := x"001f";
    tmp(41485) := x"001f";
    tmp(41486) := x"001f";
    tmp(41487) := x"001f";
    tmp(41488) := x"001f";
    tmp(41489) := x"001f";
    tmp(41490) := x"001f";
    tmp(41491) := x"001f";
    tmp(41492) := x"001f";
    tmp(41493) := x"001f";
    tmp(41494) := x"001f";
    tmp(41495) := x"001f";
    tmp(41496) := x"001f";
    tmp(41497) := x"001f";
    tmp(41498) := x"001f";
    tmp(41499) := x"001f";
    tmp(41500) := x"001f";
    tmp(41501) := x"001f";
    tmp(41502) := x"001f";
    tmp(41503) := x"001f";
    tmp(41504) := x"001f";
    tmp(41505) := x"001f";
    tmp(41506) := x"001f";
    tmp(41507) := x"001f";
    tmp(41508) := x"001f";
    tmp(41509) := x"001f";
    tmp(41510) := x"001f";
    tmp(41511) := x"001f";
    tmp(41512) := x"001f";
    tmp(41513) := x"001f";
    tmp(41514) := x"001f";
    tmp(41515) := x"001f";
    tmp(41516) := x"001f";
    tmp(41517) := x"1061";
    tmp(41518) := x"1061";
    tmp(41519) := x"1061";
    tmp(41520) := x"0000";
    tmp(41521) := x"0860";
    tmp(41522) := x"0860";
    tmp(41523) := x"0860";
    tmp(41524) := x"0860";
    tmp(41525) := x"0860";
    tmp(41526) := x"0860";
    tmp(41527) := x"0840";
    tmp(41528) := x"0840";
    tmp(41529) := x"0860";
    tmp(41530) := x"0840";
    tmp(41531) := x"0840";
    tmp(41532) := x"0860";
    tmp(41533) := x"0860";
    tmp(41534) := x"0860";
    tmp(41535) := x"0860";
    tmp(41536) := x"0860";
    tmp(41537) := x"0860";
    tmp(41538) := x"0860";
    tmp(41539) := x"0880";
    tmp(41540) := x"0880";
    tmp(41541) := x"0880";
    tmp(41542) := x"0880";
    tmp(41543) := x"08a0";
    tmp(41544) := x"08a0";
    tmp(41545) := x"08a0";
    tmp(41546) := x"08c0";
    tmp(41547) := x"08c0";
    tmp(41548) := x"08c0";
    tmp(41549) := x"08c0";
    tmp(41550) := x"08e0";
    tmp(41551) := x"08e0";
    tmp(41552) := x"08e0";
    tmp(41553) := x"0900";
    tmp(41554) := x"0900";
    tmp(41555) := x"0900";
    tmp(41556) := x"0900";
    tmp(41557) := x"0900";
    tmp(41558) := x"0920";
    tmp(41559) := x"0920";
    tmp(41560) := x"0920";
    tmp(41561) := x"0920";
    tmp(41562) := x"1140";
    tmp(41563) := x"1140";
    tmp(41564) := x"1140";
    tmp(41565) := x"1120";
    tmp(41566) := x"1140";
    tmp(41567) := x"1120";
    tmp(41568) := x"0920";
    tmp(41569) := x"1140";
    tmp(41570) := x"1140";
    tmp(41571) := x"1160";
    tmp(41572) := x"1161";
    tmp(41573) := x"1161";
    tmp(41574) := x"1161";
    tmp(41575) := x"1141";
    tmp(41576) := x"1140";
    tmp(41577) := x"1140";
    tmp(41578) := x"1140";
    tmp(41579) := x"1120";
    tmp(41580) := x"1141";
    tmp(41581) := x"1120";
    tmp(41582) := x"1140";
    tmp(41583) := x"1140";
    tmp(41584) := x"1120";
    tmp(41585) := x"1120";
    tmp(41586) := x"0920";
    tmp(41587) := x"0920";
    tmp(41588) := x"0920";
    tmp(41589) := x"0920";
    tmp(41590) := x"0920";
    tmp(41591) := x"0920";
    tmp(41592) := x"0920";
    tmp(41593) := x"0920";
    tmp(41594) := x"0940";
    tmp(41595) := x"0920";
    tmp(41596) := x"0920";
    tmp(41597) := x"0920";
    tmp(41598) := x"0920";
    tmp(41599) := x"0920";
    tmp(41600) := x"0920";
    tmp(41601) := x"0900";
    tmp(41602) := x"0900";
    tmp(41603) := x"0920";
    tmp(41604) := x"0900";
    tmp(41605) := x"0920";
    tmp(41606) := x"0900";
    tmp(41607) := x"0900";
    tmp(41608) := x"0900";
    tmp(41609) := x"0900";
    tmp(41610) := x"0900";
    tmp(41611) := x"0900";
    tmp(41612) := x"0900";
    tmp(41613) := x"0920";
    tmp(41614) := x"0900";
    tmp(41615) := x"0900";
    tmp(41616) := x"0900";
    tmp(41617) := x"0900";
    tmp(41618) := x"0920";
    tmp(41619) := x"0900";
    tmp(41620) := x"0900";
    tmp(41621) := x"0900";
    tmp(41622) := x"0900";
    tmp(41623) := x"0900";
    tmp(41624) := x"0900";
    tmp(41625) := x"0900";
    tmp(41626) := x"0900";
    tmp(41627) := x"08e0";
    tmp(41628) := x"08e0";
    tmp(41629) := x"08e0";
    tmp(41630) := x"08e0";
    tmp(41631) := x"08c0";
    tmp(41632) := x"08c0";
    tmp(41633) := x"08c0";
    tmp(41634) := x"08c0";
    tmp(41635) := x"08a0";
    tmp(41636) := x"08a0";
    tmp(41637) := x"08a0";
    tmp(41638) := x"08a0";
    tmp(41639) := x"08a0";
    tmp(41640) := x"0880";
    tmp(41641) := x"0880";
    tmp(41642) := x"2121";
    tmp(41643) := x"6ae5";
    tmp(41644) := x"b409";
    tmp(41645) := x"b389";
    tmp(41646) := x"aac7";
    tmp(41647) := x"a287";
    tmp(41648) := x"aa87";
    tmp(41649) := x"aaa7";
    tmp(41650) := x"b309";
    tmp(41651) := x"e46d";
    tmp(41652) := x"ecce";
    tmp(41653) := x"e44d";
    tmp(41654) := x"eccf";
    tmp(41655) := x"fdf2";
    tmp(41656) := x"fdb2";
    tmp(41657) := x"fd51";
    tmp(41658) := x"f48d";
    tmp(41659) := x"ec4c";
    tmp(41660) := x"ec8d";
    tmp(41661) := x"f4ce";
    tmp(41662) := x"ec8d";
    tmp(41663) := x"fcce";
    tmp(41664) := x"fcad";
    tmp(41665) := x"fd0e";
    tmp(41666) := x"f4ee";
    tmp(41667) := x"fd2f";
    tmp(41668) := x"fd10";
    tmp(41669) := x"fdb2";
    tmp(41670) := x"fdf4";
    tmp(41671) := x"fdf4";
    tmp(41672) := x"fe36";
    tmp(41673) := x"fdf5";
    tmp(41674) := x"f5f4";
    tmp(41675) := x"d48e";
    tmp(41676) := x"9205";
    tmp(41677) := x"3040";
    tmp(41678) := x"1000";
    tmp(41679) := x"1800";
    tmp(41680) := x"1800";
    tmp(41681) := x"1800";
    tmp(41682) := x"2800";
    tmp(41683) := x"3000";
    tmp(41684) := x"3000";
    tmp(41685) := x"3000";
    tmp(41686) := x"4000";
    tmp(41687) := x"5000";
    tmp(41688) := x"6820";
    tmp(41689) := x"8820";
    tmp(41690) := x"a841";
    tmp(41691) := x"c861";
    tmp(41692) := x"d081";
    tmp(41693) := x"6881";
    tmp(41694) := x"1840";
    tmp(41695) := x"1040";
    tmp(41696) := x"1040";
    tmp(41697) := x"0840";
    tmp(41698) := x"1060";
    tmp(41699) := x"1040";
    tmp(41700) := x"1040";
    tmp(41701) := x"1061";
    tmp(41702) := x"1060";
    tmp(41703) := x"1040";
    tmp(41704) := x"1040";
    tmp(41705) := x"1040";
    tmp(41706) := x"1040";
    tmp(41707) := x"0840";
    tmp(41708) := x"0840";
    tmp(41709) := x"0840";
    tmp(41710) := x"0840";
    tmp(41711) := x"0840";
    tmp(41712) := x"0840";
    tmp(41713) := x"0840";
    tmp(41714) := x"0840";
    tmp(41715) := x"0840";
    tmp(41716) := x"0840";
    tmp(41717) := x"001f";
    tmp(41718) := x"001f";
    tmp(41719) := x"001f";
    tmp(41720) := x"001f";
    tmp(41721) := x"001f";
    tmp(41722) := x"001f";
    tmp(41723) := x"001f";
    tmp(41724) := x"001f";
    tmp(41725) := x"001f";
    tmp(41726) := x"001f";
    tmp(41727) := x"001f";
    tmp(41728) := x"001f";
    tmp(41729) := x"001f";
    tmp(41730) := x"001f";
    tmp(41731) := x"001f";
    tmp(41732) := x"001f";
    tmp(41733) := x"001f";
    tmp(41734) := x"001f";
    tmp(41735) := x"001f";
    tmp(41736) := x"001f";
    tmp(41737) := x"001f";
    tmp(41738) := x"001f";
    tmp(41739) := x"001f";
    tmp(41740) := x"001f";
    tmp(41741) := x"001f";
    tmp(41742) := x"001f";
    tmp(41743) := x"001f";
    tmp(41744) := x"001f";
    tmp(41745) := x"001f";
    tmp(41746) := x"001f";
    tmp(41747) := x"001f";
    tmp(41748) := x"001f";
    tmp(41749) := x"001f";
    tmp(41750) := x"001f";
    tmp(41751) := x"001f";
    tmp(41752) := x"001f";
    tmp(41753) := x"001f";
    tmp(41754) := x"001f";
    tmp(41755) := x"001f";
    tmp(41756) := x"001f";
    tmp(41757) := x"1061";
    tmp(41758) := x"1061";
    tmp(41759) := x"1061";
    tmp(41760) := x"0000";
    tmp(41761) := x"0860";
    tmp(41762) := x"0860";
    tmp(41763) := x"0860";
    tmp(41764) := x"0860";
    tmp(41765) := x"0860";
    tmp(41766) := x"0860";
    tmp(41767) := x"0840";
    tmp(41768) := x"0840";
    tmp(41769) := x"0840";
    tmp(41770) := x"0860";
    tmp(41771) := x"0840";
    tmp(41772) := x"0840";
    tmp(41773) := x"0840";
    tmp(41774) := x"0860";
    tmp(41775) := x"0860";
    tmp(41776) := x"0860";
    tmp(41777) := x"0860";
    tmp(41778) := x"0860";
    tmp(41779) := x"0860";
    tmp(41780) := x"0860";
    tmp(41781) := x"0880";
    tmp(41782) := x"0880";
    tmp(41783) := x"0880";
    tmp(41784) := x"08a0";
    tmp(41785) := x"08a0";
    tmp(41786) := x"08a0";
    tmp(41787) := x"08c0";
    tmp(41788) := x"08c0";
    tmp(41789) := x"08c0";
    tmp(41790) := x"08c0";
    tmp(41791) := x"08e0";
    tmp(41792) := x"08e0";
    tmp(41793) := x"08e0";
    tmp(41794) := x"08e0";
    tmp(41795) := x"08e0";
    tmp(41796) := x"0900";
    tmp(41797) := x"0900";
    tmp(41798) := x"0920";
    tmp(41799) := x"0920";
    tmp(41800) := x"0920";
    tmp(41801) := x"0920";
    tmp(41802) := x"0920";
    tmp(41803) := x"0940";
    tmp(41804) := x"0940";
    tmp(41805) := x"0920";
    tmp(41806) := x"0920";
    tmp(41807) := x"0920";
    tmp(41808) := x"0920";
    tmp(41809) := x"0920";
    tmp(41810) := x"1140";
    tmp(41811) := x"1140";
    tmp(41812) := x"1140";
    tmp(41813) := x"1140";
    tmp(41814) := x"1161";
    tmp(41815) := x"1141";
    tmp(41816) := x"1140";
    tmp(41817) := x"1140";
    tmp(41818) := x"1120";
    tmp(41819) := x"1120";
    tmp(41820) := x"1120";
    tmp(41821) := x"1120";
    tmp(41822) := x"1140";
    tmp(41823) := x"1140";
    tmp(41824) := x"1120";
    tmp(41825) := x"1120";
    tmp(41826) := x"0920";
    tmp(41827) := x"0920";
    tmp(41828) := x"0940";
    tmp(41829) := x"0920";
    tmp(41830) := x"0920";
    tmp(41831) := x"0920";
    tmp(41832) := x"0920";
    tmp(41833) := x"0920";
    tmp(41834) := x"0920";
    tmp(41835) := x"0920";
    tmp(41836) := x"0920";
    tmp(41837) := x"0920";
    tmp(41838) := x"0920";
    tmp(41839) := x"0920";
    tmp(41840) := x"0920";
    tmp(41841) := x"0920";
    tmp(41842) := x"0900";
    tmp(41843) := x"0920";
    tmp(41844) := x"0900";
    tmp(41845) := x"0920";
    tmp(41846) := x"0900";
    tmp(41847) := x"0900";
    tmp(41848) := x"0900";
    tmp(41849) := x"0900";
    tmp(41850) := x"0900";
    tmp(41851) := x"0900";
    tmp(41852) := x"0900";
    tmp(41853) := x"0900";
    tmp(41854) := x"0900";
    tmp(41855) := x"0900";
    tmp(41856) := x"0900";
    tmp(41857) := x"0920";
    tmp(41858) := x"0920";
    tmp(41859) := x"0900";
    tmp(41860) := x"0900";
    tmp(41861) := x"0920";
    tmp(41862) := x"0900";
    tmp(41863) := x"0900";
    tmp(41864) := x"0900";
    tmp(41865) := x"0900";
    tmp(41866) := x"0900";
    tmp(41867) := x"08e0";
    tmp(41868) := x"08e0";
    tmp(41869) := x"08c0";
    tmp(41870) := x"08e0";
    tmp(41871) := x"08c0";
    tmp(41872) := x"08c0";
    tmp(41873) := x"08c0";
    tmp(41874) := x"08c0";
    tmp(41875) := x"08a0";
    tmp(41876) := x"08a0";
    tmp(41877) := x"08a0";
    tmp(41878) := x"0880";
    tmp(41879) := x"10a0";
    tmp(41880) := x"41e2";
    tmp(41881) := x"a3a7";
    tmp(41882) := x"bbe9";
    tmp(41883) := x"ab27";
    tmp(41884) := x"a286";
    tmp(41885) := x"baa7";
    tmp(41886) := x"c2c7";
    tmp(41887) := x"cb08";
    tmp(41888) := x"d328";
    tmp(41889) := x"cb08";
    tmp(41890) := x"baa7";
    tmp(41891) := x"c329";
    tmp(41892) := x"ecce";
    tmp(41893) := x"ec6d";
    tmp(41894) := x"e40d";
    tmp(41895) := x"f4cf";
    tmp(41896) := x"fd71";
    tmp(41897) := x"fd30";
    tmp(41898) := x"f48d";
    tmp(41899) := x"fd2f";
    tmp(41900) := x"fd91";
    tmp(41901) := x"fd10";
    tmp(41902) := x"fd50";
    tmp(41903) := x"fcee";
    tmp(41904) := x"fc6d";
    tmp(41905) := x"fc8d";
    tmp(41906) := x"fcad";
    tmp(41907) := x"fcef";
    tmp(41908) := x"fd71";
    tmp(41909) := x"fd31";
    tmp(41910) := x"fdb2";
    tmp(41911) := x"fdd3";
    tmp(41912) := x"fdf4";
    tmp(41913) := x"fd93";
    tmp(41914) := x"f4b1";
    tmp(41915) := x"cb4b";
    tmp(41916) := x"50c2";
    tmp(41917) := x"2020";
    tmp(41918) := x"1800";
    tmp(41919) := x"1000";
    tmp(41920) := x"1000";
    tmp(41921) := x"1000";
    tmp(41922) := x"2000";
    tmp(41923) := x"2800";
    tmp(41924) := x"2800";
    tmp(41925) := x"3000";
    tmp(41926) := x"3800";
    tmp(41927) := x"5000";
    tmp(41928) := x"6000";
    tmp(41929) := x"7820";
    tmp(41930) := x"8820";
    tmp(41931) := x"9820";
    tmp(41932) := x"a841";
    tmp(41933) := x"c881";
    tmp(41934) := x"6081";
    tmp(41935) := x"1840";
    tmp(41936) := x"1040";
    tmp(41937) := x"1040";
    tmp(41938) := x"0840";
    tmp(41939) := x"1040";
    tmp(41940) := x"1040";
    tmp(41941) := x"1040";
    tmp(41942) := x"1040";
    tmp(41943) := x"1040";
    tmp(41944) := x"1060";
    tmp(41945) := x"1040";
    tmp(41946) := x"0840";
    tmp(41947) := x"0840";
    tmp(41948) := x"0840";
    tmp(41949) := x"0840";
    tmp(41950) := x"0840";
    tmp(41951) := x"0840";
    tmp(41952) := x"0840";
    tmp(41953) := x"0840";
    tmp(41954) := x"0840";
    tmp(41955) := x"0840";
    tmp(41956) := x"0840";
    tmp(41957) := x"001f";
    tmp(41958) := x"001f";
    tmp(41959) := x"001f";
    tmp(41960) := x"001f";
    tmp(41961) := x"001f";
    tmp(41962) := x"001f";
    tmp(41963) := x"001f";
    tmp(41964) := x"001f";
    tmp(41965) := x"001f";
    tmp(41966) := x"001f";
    tmp(41967) := x"001f";
    tmp(41968) := x"001f";
    tmp(41969) := x"001f";
    tmp(41970) := x"001f";
    tmp(41971) := x"001f";
    tmp(41972) := x"001f";
    tmp(41973) := x"001f";
    tmp(41974) := x"001f";
    tmp(41975) := x"001f";
    tmp(41976) := x"001f";
    tmp(41977) := x"001f";
    tmp(41978) := x"001f";
    tmp(41979) := x"001f";
    tmp(41980) := x"001f";
    tmp(41981) := x"001f";
    tmp(41982) := x"001f";
    tmp(41983) := x"001f";
    tmp(41984) := x"001f";
    tmp(41985) := x"001f";
    tmp(41986) := x"001f";
    tmp(41987) := x"001f";
    tmp(41988) := x"001f";
    tmp(41989) := x"001f";
    tmp(41990) := x"001f";
    tmp(41991) := x"001f";
    tmp(41992) := x"001f";
    tmp(41993) := x"001f";
    tmp(41994) := x"001f";
    tmp(41995) := x"001f";
    tmp(41996) := x"001f";
    tmp(41997) := x"1061";
    tmp(41998) := x"1061";
    tmp(41999) := x"1061";
    tmp(42000) := x"0000";
    tmp(42001) := x"0860";
    tmp(42002) := x"0860";
    tmp(42003) := x"0860";
    tmp(42004) := x"0860";
    tmp(42005) := x"0860";
    tmp(42006) := x"0860";
    tmp(42007) := x"0840";
    tmp(42008) := x"0840";
    tmp(42009) := x"0840";
    tmp(42010) := x"0840";
    tmp(42011) := x"0840";
    tmp(42012) := x"0840";
    tmp(42013) := x"0840";
    tmp(42014) := x"0840";
    tmp(42015) := x"0840";
    tmp(42016) := x"0860";
    tmp(42017) := x"0860";
    tmp(42018) := x"0860";
    tmp(42019) := x"0860";
    tmp(42020) := x"0860";
    tmp(42021) := x"0860";
    tmp(42022) := x"0860";
    tmp(42023) := x"0880";
    tmp(42024) := x"0880";
    tmp(42025) := x"08a0";
    tmp(42026) := x"08a0";
    tmp(42027) := x"08a0";
    tmp(42028) := x"08c0";
    tmp(42029) := x"08c0";
    tmp(42030) := x"08c0";
    tmp(42031) := x"08c0";
    tmp(42032) := x"08e0";
    tmp(42033) := x"08e0";
    tmp(42034) := x"08e0";
    tmp(42035) := x"08e0";
    tmp(42036) := x"08e0";
    tmp(42037) := x"0900";
    tmp(42038) := x"0900";
    tmp(42039) := x"0900";
    tmp(42040) := x"0900";
    tmp(42041) := x"0920";
    tmp(42042) := x"0920";
    tmp(42043) := x"0920";
    tmp(42044) := x"0920";
    tmp(42045) := x"0920";
    tmp(42046) := x"0920";
    tmp(42047) := x"0920";
    tmp(42048) := x"0920";
    tmp(42049) := x"0920";
    tmp(42050) := x"0920";
    tmp(42051) := x"1140";
    tmp(42052) := x"1140";
    tmp(42053) := x"1140";
    tmp(42054) := x"1140";
    tmp(42055) := x"1140";
    tmp(42056) := x"1140";
    tmp(42057) := x"1120";
    tmp(42058) := x"1120";
    tmp(42059) := x"0920";
    tmp(42060) := x"1120";
    tmp(42061) := x"1120";
    tmp(42062) := x"1120";
    tmp(42063) := x"1120";
    tmp(42064) := x"1140";
    tmp(42065) := x"1140";
    tmp(42066) := x"0920";
    tmp(42067) := x"0940";
    tmp(42068) := x"0920";
    tmp(42069) := x"0920";
    tmp(42070) := x"0920";
    tmp(42071) := x"0920";
    tmp(42072) := x"0920";
    tmp(42073) := x"0920";
    tmp(42074) := x"0920";
    tmp(42075) := x"0920";
    tmp(42076) := x"0920";
    tmp(42077) := x"0920";
    tmp(42078) := x"0920";
    tmp(42079) := x"0920";
    tmp(42080) := x"0900";
    tmp(42081) := x"0900";
    tmp(42082) := x"0920";
    tmp(42083) := x"0920";
    tmp(42084) := x"0900";
    tmp(42085) := x"0900";
    tmp(42086) := x"0900";
    tmp(42087) := x"0900";
    tmp(42088) := x"0900";
    tmp(42089) := x"0900";
    tmp(42090) := x"0900";
    tmp(42091) := x"0900";
    tmp(42092) := x"0900";
    tmp(42093) := x"0900";
    tmp(42094) := x"0900";
    tmp(42095) := x"0900";
    tmp(42096) := x"0900";
    tmp(42097) := x"0920";
    tmp(42098) := x"0920";
    tmp(42099) := x"0900";
    tmp(42100) := x"0900";
    tmp(42101) := x"0900";
    tmp(42102) := x"0900";
    tmp(42103) := x"0920";
    tmp(42104) := x"0900";
    tmp(42105) := x"08e0";
    tmp(42106) := x"08e0";
    tmp(42107) := x"08e0";
    tmp(42108) := x"08e0";
    tmp(42109) := x"08e0";
    tmp(42110) := x"08c0";
    tmp(42111) := x"08c0";
    tmp(42112) := x"08c0";
    tmp(42113) := x"08c0";
    tmp(42114) := x"08a0";
    tmp(42115) := x"08a0";
    tmp(42116) := x"08a0";
    tmp(42117) := x"0880";
    tmp(42118) := x"3181";
    tmp(42119) := x"82e5";
    tmp(42120) := x"ab48";
    tmp(42121) := x"a2a7";
    tmp(42122) := x"aaa7";
    tmp(42123) := x"bac7";
    tmp(42124) := x"c308";
    tmp(42125) := x"d348";
    tmp(42126) := x"cb28";
    tmp(42127) := x"db49";
    tmp(42128) := x"d349";
    tmp(42129) := x"c308";
    tmp(42130) := x"cac8";
    tmp(42131) := x"b2a7";
    tmp(42132) := x"ec8d";
    tmp(42133) := x"ec6e";
    tmp(42134) := x"dbac";
    tmp(42135) := x"e3ed";
    tmp(42136) := x"fcf0";
    tmp(42137) := x"ec6e";
    tmp(42138) := x"fcae";
    tmp(42139) := x"f48e";
    tmp(42140) := x"fcaf";
    tmp(42141) := x"fc8e";
    tmp(42142) := x"fc8e";
    tmp(42143) := x"fcae";
    tmp(42144) := x"fcef";
    tmp(42145) := x"fcef";
    tmp(42146) := x"fcae";
    tmp(42147) := x"fd31";
    tmp(42148) := x"fd31";
    tmp(42149) := x"fcf0";
    tmp(42150) := x"fd31";
    tmp(42151) := x"fd51";
    tmp(42152) := x"fdb3";
    tmp(42153) := x"f532";
    tmp(42154) := x"e44f";
    tmp(42155) := x"bac8";
    tmp(42156) := x"58c2";
    tmp(42157) := x"1800";
    tmp(42158) := x"1000";
    tmp(42159) := x"1000";
    tmp(42160) := x"1000";
    tmp(42161) := x"1000";
    tmp(42162) := x"1800";
    tmp(42163) := x"1800";
    tmp(42164) := x"2800";
    tmp(42165) := x"3800";
    tmp(42166) := x"4000";
    tmp(42167) := x"4000";
    tmp(42168) := x"4800";
    tmp(42169) := x"5000";
    tmp(42170) := x"6000";
    tmp(42171) := x"8020";
    tmp(42172) := x"8820";
    tmp(42173) := x"b021";
    tmp(42174) := x"e081";
    tmp(42175) := x"6881";
    tmp(42176) := x"1840";
    tmp(42177) := x"1040";
    tmp(42178) := x"1040";
    tmp(42179) := x"1040";
    tmp(42180) := x"1040";
    tmp(42181) := x"1040";
    tmp(42182) := x"0840";
    tmp(42183) := x"1040";
    tmp(42184) := x"1040";
    tmp(42185) := x"0840";
    tmp(42186) := x"0840";
    tmp(42187) := x"0840";
    tmp(42188) := x"0840";
    tmp(42189) := x"0840";
    tmp(42190) := x"0840";
    tmp(42191) := x"0840";
    tmp(42192) := x"0840";
    tmp(42193) := x"0840";
    tmp(42194) := x"0840";
    tmp(42195) := x"0840";
    tmp(42196) := x"0840";
    tmp(42197) := x"001f";
    tmp(42198) := x"001f";
    tmp(42199) := x"001f";
    tmp(42200) := x"001f";
    tmp(42201) := x"001f";
    tmp(42202) := x"001f";
    tmp(42203) := x"001f";
    tmp(42204) := x"001f";
    tmp(42205) := x"001f";
    tmp(42206) := x"001f";
    tmp(42207) := x"001f";
    tmp(42208) := x"001f";
    tmp(42209) := x"001f";
    tmp(42210) := x"001f";
    tmp(42211) := x"001f";
    tmp(42212) := x"001f";
    tmp(42213) := x"001f";
    tmp(42214) := x"001f";
    tmp(42215) := x"001f";
    tmp(42216) := x"001f";
    tmp(42217) := x"001f";
    tmp(42218) := x"001f";
    tmp(42219) := x"001f";
    tmp(42220) := x"001f";
    tmp(42221) := x"001f";
    tmp(42222) := x"001f";
    tmp(42223) := x"001f";
    tmp(42224) := x"001f";
    tmp(42225) := x"001f";
    tmp(42226) := x"001f";
    tmp(42227) := x"001f";
    tmp(42228) := x"001f";
    tmp(42229) := x"001f";
    tmp(42230) := x"001f";
    tmp(42231) := x"001f";
    tmp(42232) := x"001f";
    tmp(42233) := x"001f";
    tmp(42234) := x"001f";
    tmp(42235) := x"001f";
    tmp(42236) := x"001f";
    tmp(42237) := x"1061";
    tmp(42238) := x"1061";
    tmp(42239) := x"1061";
    tmp(42240) := x"0000";
    tmp(42241) := x"0880";
    tmp(42242) := x"0880";
    tmp(42243) := x"0860";
    tmp(42244) := x"0860";
    tmp(42245) := x"0860";
    tmp(42246) := x"0860";
    tmp(42247) := x"0860";
    tmp(42248) := x"0860";
    tmp(42249) := x"0860";
    tmp(42250) := x"0840";
    tmp(42251) := x"0840";
    tmp(42252) := x"0840";
    tmp(42253) := x"0840";
    tmp(42254) := x"0840";
    tmp(42255) := x"0840";
    tmp(42256) := x"0840";
    tmp(42257) := x"0860";
    tmp(42258) := x"0860";
    tmp(42259) := x"0860";
    tmp(42260) := x"0860";
    tmp(42261) := x"0860";
    tmp(42262) := x"0860";
    tmp(42263) := x"0860";
    tmp(42264) := x"0880";
    tmp(42265) := x"0880";
    tmp(42266) := x"08a0";
    tmp(42267) := x"08a0";
    tmp(42268) := x"08a0";
    tmp(42269) := x"08c0";
    tmp(42270) := x"08c0";
    tmp(42271) := x"08c0";
    tmp(42272) := x"08e0";
    tmp(42273) := x"08e0";
    tmp(42274) := x"08e0";
    tmp(42275) := x"08e0";
    tmp(42276) := x"08e0";
    tmp(42277) := x"08e0";
    tmp(42278) := x"0900";
    tmp(42279) := x"0900";
    tmp(42280) := x"0900";
    tmp(42281) := x"0900";
    tmp(42282) := x"0920";
    tmp(42283) := x"0920";
    tmp(42284) := x"0920";
    tmp(42285) := x"0920";
    tmp(42286) := x"0920";
    tmp(42287) := x"0900";
    tmp(42288) := x"0920";
    tmp(42289) := x"0900";
    tmp(42290) := x"0920";
    tmp(42291) := x"0920";
    tmp(42292) := x"1140";
    tmp(42293) := x"1140";
    tmp(42294) := x"1140";
    tmp(42295) := x"1120";
    tmp(42296) := x"1120";
    tmp(42297) := x"1120";
    tmp(42298) := x"0920";
    tmp(42299) := x"1120";
    tmp(42300) := x"1120";
    tmp(42301) := x"0920";
    tmp(42302) := x"0920";
    tmp(42303) := x"1120";
    tmp(42304) := x"0920";
    tmp(42305) := x"0920";
    tmp(42306) := x"0920";
    tmp(42307) := x"1140";
    tmp(42308) := x"0940";
    tmp(42309) := x"0920";
    tmp(42310) := x"0920";
    tmp(42311) := x"0920";
    tmp(42312) := x"0920";
    tmp(42313) := x"0920";
    tmp(42314) := x"0920";
    tmp(42315) := x"0920";
    tmp(42316) := x"0920";
    tmp(42317) := x"0920";
    tmp(42318) := x"0920";
    tmp(42319) := x"0920";
    tmp(42320) := x"0920";
    tmp(42321) := x"0920";
    tmp(42322) := x"0900";
    tmp(42323) := x"0900";
    tmp(42324) := x"0900";
    tmp(42325) := x"0900";
    tmp(42326) := x"0900";
    tmp(42327) := x"0900";
    tmp(42328) := x"0900";
    tmp(42329) := x"0900";
    tmp(42330) := x"0900";
    tmp(42331) := x"0900";
    tmp(42332) := x"0900";
    tmp(42333) := x"0900";
    tmp(42334) := x"0900";
    tmp(42335) := x"0920";
    tmp(42336) := x"0920";
    tmp(42337) := x"0920";
    tmp(42338) := x"0920";
    tmp(42339) := x"0900";
    tmp(42340) := x"0920";
    tmp(42341) := x"0900";
    tmp(42342) := x"0920";
    tmp(42343) := x"0900";
    tmp(42344) := x"0900";
    tmp(42345) := x"0900";
    tmp(42346) := x"0900";
    tmp(42347) := x"08e0";
    tmp(42348) := x"08e0";
    tmp(42349) := x"08e0";
    tmp(42350) := x"08c0";
    tmp(42351) := x"08c0";
    tmp(42352) := x"08a0";
    tmp(42353) := x"08a0";
    tmp(42354) := x"08a0";
    tmp(42355) := x"08a0";
    tmp(42356) := x"18e0";
    tmp(42357) := x"5a03";
    tmp(42358) := x"7a04";
    tmp(42359) := x"8a45";
    tmp(42360) := x"a287";
    tmp(42361) := x"bb08";
    tmp(42362) := x"bb08";
    tmp(42363) := x"c349";
    tmp(42364) := x"c349";
    tmp(42365) := x"c328";
    tmp(42366) := x"cb29";
    tmp(42367) := x"cb29";
    tmp(42368) := x"cb09";
    tmp(42369) := x"cb09";
    tmp(42370) := x"c2c8";
    tmp(42371) := x"bae8";
    tmp(42372) := x"ec2d";
    tmp(42373) := x"cb8b";
    tmp(42374) := x"cb6a";
    tmp(42375) := x"dbab";
    tmp(42376) := x"dbab";
    tmp(42377) := x"dbab";
    tmp(42378) := x"ebec";
    tmp(42379) := x"f42d";
    tmp(42380) := x"ec0d";
    tmp(42381) := x"f46e";
    tmp(42382) := x"fc8e";
    tmp(42383) := x"f46e";
    tmp(42384) := x"fcaf";
    tmp(42385) := x"fccf";
    tmp(42386) := x"fd31";
    tmp(42387) := x"fcf1";
    tmp(42388) := x"fcf2";
    tmp(42389) := x"fd52";
    tmp(42390) := x"fd32";
    tmp(42391) := x"fd12";
    tmp(42392) := x"f511";
    tmp(42393) := x"ec70";
    tmp(42394) := x"dbee";
    tmp(42395) := x"b2a8";
    tmp(42396) := x"60e2";
    tmp(42397) := x"1800";
    tmp(42398) := x"0800";
    tmp(42399) := x"1000";
    tmp(42400) := x"1000";
    tmp(42401) := x"1000";
    tmp(42402) := x"1000";
    tmp(42403) := x"1000";
    tmp(42404) := x"2000";
    tmp(42405) := x"3000";
    tmp(42406) := x"3800";
    tmp(42407) := x"3800";
    tmp(42408) := x"3800";
    tmp(42409) := x"4000";
    tmp(42410) := x"5000";
    tmp(42411) := x"7800";
    tmp(42412) := x"9020";
    tmp(42413) := x"9820";
    tmp(42414) := x"c021";
    tmp(42415) := x"d061";
    tmp(42416) := x"3861";
    tmp(42417) := x"1040";
    tmp(42418) := x"1040";
    tmp(42419) := x"1040";
    tmp(42420) := x"0840";
    tmp(42421) := x"1040";
    tmp(42422) := x"1040";
    tmp(42423) := x"1040";
    tmp(42424) := x"0840";
    tmp(42425) := x"0840";
    tmp(42426) := x"0840";
    tmp(42427) := x"0840";
    tmp(42428) := x"0840";
    tmp(42429) := x"0840";
    tmp(42430) := x"0840";
    tmp(42431) := x"0840";
    tmp(42432) := x"0840";
    tmp(42433) := x"0840";
    tmp(42434) := x"0840";
    tmp(42435) := x"0840";
    tmp(42436) := x"0840";
    tmp(42437) := x"001f";
    tmp(42438) := x"001f";
    tmp(42439) := x"001f";
    tmp(42440) := x"001f";
    tmp(42441) := x"001f";
    tmp(42442) := x"001f";
    tmp(42443) := x"001f";
    tmp(42444) := x"001f";
    tmp(42445) := x"001f";
    tmp(42446) := x"001f";
    tmp(42447) := x"001f";
    tmp(42448) := x"001f";
    tmp(42449) := x"001f";
    tmp(42450) := x"001f";
    tmp(42451) := x"001f";
    tmp(42452) := x"001f";
    tmp(42453) := x"001f";
    tmp(42454) := x"001f";
    tmp(42455) := x"001f";
    tmp(42456) := x"001f";
    tmp(42457) := x"001f";
    tmp(42458) := x"001f";
    tmp(42459) := x"001f";
    tmp(42460) := x"001f";
    tmp(42461) := x"001f";
    tmp(42462) := x"001f";
    tmp(42463) := x"001f";
    tmp(42464) := x"001f";
    tmp(42465) := x"001f";
    tmp(42466) := x"001f";
    tmp(42467) := x"001f";
    tmp(42468) := x"001f";
    tmp(42469) := x"001f";
    tmp(42470) := x"001f";
    tmp(42471) := x"001f";
    tmp(42472) := x"001f";
    tmp(42473) := x"001f";
    tmp(42474) := x"001f";
    tmp(42475) := x"001f";
    tmp(42476) := x"001f";
    tmp(42477) := x"1061";
    tmp(42478) := x"1061";
    tmp(42479) := x"1061";
    tmp(42480) := x"0000";
    tmp(42481) := x"0880";
    tmp(42482) := x"0880";
    tmp(42483) := x"0860";
    tmp(42484) := x"0880";
    tmp(42485) := x"0860";
    tmp(42486) := x"0860";
    tmp(42487) := x"0860";
    tmp(42488) := x"0860";
    tmp(42489) := x"0860";
    tmp(42490) := x"0860";
    tmp(42491) := x"0840";
    tmp(42492) := x"0840";
    tmp(42493) := x"0840";
    tmp(42494) := x"0840";
    tmp(42495) := x"0840";
    tmp(42496) := x"0840";
    tmp(42497) := x"0840";
    tmp(42498) := x"0840";
    tmp(42499) := x"0840";
    tmp(42500) := x"0840";
    tmp(42501) := x"0860";
    tmp(42502) := x"0860";
    tmp(42503) := x"0860";
    tmp(42504) := x"0860";
    tmp(42505) := x"0860";
    tmp(42506) := x"0880";
    tmp(42507) := x"08a0";
    tmp(42508) := x"08a0";
    tmp(42509) := x"08a0";
    tmp(42510) := x"08c0";
    tmp(42511) := x"08c0";
    tmp(42512) := x"08c0";
    tmp(42513) := x"08c0";
    tmp(42514) := x"08c0";
    tmp(42515) := x"08e0";
    tmp(42516) := x"08e0";
    tmp(42517) := x"08e0";
    tmp(42518) := x"08e0";
    tmp(42519) := x"0900";
    tmp(42520) := x"0900";
    tmp(42521) := x"0900";
    tmp(42522) := x"0900";
    tmp(42523) := x"0920";
    tmp(42524) := x"0920";
    tmp(42525) := x"0920";
    tmp(42526) := x"0920";
    tmp(42527) := x"0900";
    tmp(42528) := x"0900";
    tmp(42529) := x"0920";
    tmp(42530) := x"0920";
    tmp(42531) := x"0920";
    tmp(42532) := x"0920";
    tmp(42533) := x"1140";
    tmp(42534) := x"1120";
    tmp(42535) := x"1140";
    tmp(42536) := x"1140";
    tmp(42537) := x"1120";
    tmp(42538) := x"1140";
    tmp(42539) := x"1120";
    tmp(42540) := x"1120";
    tmp(42541) := x"0920";
    tmp(42542) := x"0920";
    tmp(42543) := x"0920";
    tmp(42544) := x"0920";
    tmp(42545) := x"0920";
    tmp(42546) := x"0920";
    tmp(42547) := x"0920";
    tmp(42548) := x"0920";
    tmp(42549) := x"0940";
    tmp(42550) := x"0940";
    tmp(42551) := x"0920";
    tmp(42552) := x"0920";
    tmp(42553) := x"0900";
    tmp(42554) := x"0900";
    tmp(42555) := x"0900";
    tmp(42556) := x"0920";
    tmp(42557) := x"0900";
    tmp(42558) := x"0900";
    tmp(42559) := x"0900";
    tmp(42560) := x"0900";
    tmp(42561) := x"0900";
    tmp(42562) := x"0900";
    tmp(42563) := x"0900";
    tmp(42564) := x"0900";
    tmp(42565) := x"0900";
    tmp(42566) := x"0900";
    tmp(42567) := x"0900";
    tmp(42568) := x"0900";
    tmp(42569) := x"0900";
    tmp(42570) := x"0900";
    tmp(42571) := x"0900";
    tmp(42572) := x"0900";
    tmp(42573) := x"0900";
    tmp(42574) := x"0920";
    tmp(42575) := x"0920";
    tmp(42576) := x"0920";
    tmp(42577) := x"0920";
    tmp(42578) := x"0920";
    tmp(42579) := x"0900";
    tmp(42580) := x"0920";
    tmp(42581) := x"0920";
    tmp(42582) := x"0900";
    tmp(42583) := x"0900";
    tmp(42584) := x"0900";
    tmp(42585) := x"0900";
    tmp(42586) := x"0900";
    tmp(42587) := x"08e0";
    tmp(42588) := x"08e0";
    tmp(42589) := x"08e0";
    tmp(42590) := x"08c0";
    tmp(42591) := x"08c0";
    tmp(42592) := x"08a0";
    tmp(42593) := x"08a0";
    tmp(42594) := x"10a0";
    tmp(42595) := x"3981";
    tmp(42596) := x"7a44";
    tmp(42597) := x"9a86";
    tmp(42598) := x"a286";
    tmp(42599) := x"a287";
    tmp(42600) := x"bb09";
    tmp(42601) := x"bb29";
    tmp(42602) := x"cb6a";
    tmp(42603) := x"cb6b";
    tmp(42604) := x"cb6a";
    tmp(42605) := x"cb6a";
    tmp(42606) := x"cb29";
    tmp(42607) := x"cb09";
    tmp(42608) := x"cb09";
    tmp(42609) := x"cb09";
    tmp(42610) := x"baa8";
    tmp(42611) := x"c32a";
    tmp(42612) := x"dbcc";
    tmp(42613) := x"d38b";
    tmp(42614) := x"dbcc";
    tmp(42615) := x"dbab";
    tmp(42616) := x"cb4a";
    tmp(42617) := x"e3ab";
    tmp(42618) := x"ec0c";
    tmp(42619) := x"e3cc";
    tmp(42620) := x"ec0d";
    tmp(42621) := x"fcaf";
    tmp(42622) := x"fc8f";
    tmp(42623) := x"fcaf";
    tmp(42624) := x"fccf";
    tmp(42625) := x"fcf0";
    tmp(42626) := x"fcf1";
    tmp(42627) := x"fcf1";
    tmp(42628) := x"fcd1";
    tmp(42629) := x"fd33";
    tmp(42630) := x"fcf3";
    tmp(42631) := x"f491";
    tmp(42632) := x"f4d2";
    tmp(42633) := x"ecd2";
    tmp(42634) := x"dbee";
    tmp(42635) := x"aa88";
    tmp(42636) := x"58c2";
    tmp(42637) := x"1800";
    tmp(42638) := x"0800";
    tmp(42639) := x"0800";
    tmp(42640) := x"0800";
    tmp(42641) := x"1000";
    tmp(42642) := x"1000";
    tmp(42643) := x"1000";
    tmp(42644) := x"2000";
    tmp(42645) := x"3000";
    tmp(42646) := x"3800";
    tmp(42647) := x"3000";
    tmp(42648) := x"2800";
    tmp(42649) := x"3800";
    tmp(42650) := x"5000";
    tmp(42651) := x"6800";
    tmp(42652) := x"7800";
    tmp(42653) := x"7800";
    tmp(42654) := x"9020";
    tmp(42655) := x"c041";
    tmp(42656) := x"8061";
    tmp(42657) := x"1840";
    tmp(42658) := x"1040";
    tmp(42659) := x"1040";
    tmp(42660) := x"1040";
    tmp(42661) := x"1040";
    tmp(42662) := x"0840";
    tmp(42663) := x"0840";
    tmp(42664) := x"0840";
    tmp(42665) := x"0840";
    tmp(42666) := x"0840";
    tmp(42667) := x"0840";
    tmp(42668) := x"0840";
    tmp(42669) := x"0840";
    tmp(42670) := x"0840";
    tmp(42671) := x"0840";
    tmp(42672) := x"0840";
    tmp(42673) := x"0840";
    tmp(42674) := x"0840";
    tmp(42675) := x"0840";
    tmp(42676) := x"0840";
    tmp(42677) := x"001f";
    tmp(42678) := x"001f";
    tmp(42679) := x"001f";
    tmp(42680) := x"001f";
    tmp(42681) := x"001f";
    tmp(42682) := x"001f";
    tmp(42683) := x"001f";
    tmp(42684) := x"001f";
    tmp(42685) := x"001f";
    tmp(42686) := x"001f";
    tmp(42687) := x"001f";
    tmp(42688) := x"001f";
    tmp(42689) := x"001f";
    tmp(42690) := x"001f";
    tmp(42691) := x"001f";
    tmp(42692) := x"001f";
    tmp(42693) := x"001f";
    tmp(42694) := x"001f";
    tmp(42695) := x"001f";
    tmp(42696) := x"001f";
    tmp(42697) := x"001f";
    tmp(42698) := x"001f";
    tmp(42699) := x"001f";
    tmp(42700) := x"001f";
    tmp(42701) := x"001f";
    tmp(42702) := x"001f";
    tmp(42703) := x"001f";
    tmp(42704) := x"001f";
    tmp(42705) := x"001f";
    tmp(42706) := x"001f";
    tmp(42707) := x"001f";
    tmp(42708) := x"001f";
    tmp(42709) := x"001f";
    tmp(42710) := x"001f";
    tmp(42711) := x"001f";
    tmp(42712) := x"001f";
    tmp(42713) := x"001f";
    tmp(42714) := x"001f";
    tmp(42715) := x"001f";
    tmp(42716) := x"001f";
    tmp(42717) := x"1061";
    tmp(42718) := x"1061";
    tmp(42719) := x"1061";
    tmp(42720) := x"0000";
    tmp(42721) := x"0880";
    tmp(42722) := x"0880";
    tmp(42723) := x"0880";
    tmp(42724) := x"0880";
    tmp(42725) := x"0880";
    tmp(42726) := x"0860";
    tmp(42727) := x"0860";
    tmp(42728) := x"0860";
    tmp(42729) := x"0860";
    tmp(42730) := x"0860";
    tmp(42731) := x"0840";
    tmp(42732) := x"0840";
    tmp(42733) := x"0840";
    tmp(42734) := x"0840";
    tmp(42735) := x"0840";
    tmp(42736) := x"0840";
    tmp(42737) := x"0840";
    tmp(42738) := x"0840";
    tmp(42739) := x"0840";
    tmp(42740) := x"0840";
    tmp(42741) := x"0840";
    tmp(42742) := x"0840";
    tmp(42743) := x"0860";
    tmp(42744) := x"0860";
    tmp(42745) := x"0860";
    tmp(42746) := x"0860";
    tmp(42747) := x"0880";
    tmp(42748) := x"08a0";
    tmp(42749) := x"08a0";
    tmp(42750) := x"08a0";
    tmp(42751) := x"08c0";
    tmp(42752) := x"08a0";
    tmp(42753) := x"08c0";
    tmp(42754) := x"08c0";
    tmp(42755) := x"08c0";
    tmp(42756) := x"08c0";
    tmp(42757) := x"08e0";
    tmp(42758) := x"08e0";
    tmp(42759) := x"08e0";
    tmp(42760) := x"0900";
    tmp(42761) := x"0900";
    tmp(42762) := x"0900";
    tmp(42763) := x"0920";
    tmp(42764) := x"0900";
    tmp(42765) := x"0900";
    tmp(42766) := x"0900";
    tmp(42767) := x"0920";
    tmp(42768) := x"0900";
    tmp(42769) := x"0900";
    tmp(42770) := x"0900";
    tmp(42771) := x"0900";
    tmp(42772) := x"0920";
    tmp(42773) := x"0940";
    tmp(42774) := x"0920";
    tmp(42775) := x"0920";
    tmp(42776) := x"1140";
    tmp(42777) := x"0920";
    tmp(42778) := x"0920";
    tmp(42779) := x"0920";
    tmp(42780) := x"0920";
    tmp(42781) := x"0920";
    tmp(42782) := x"0920";
    tmp(42783) := x"0920";
    tmp(42784) := x"0920";
    tmp(42785) := x"0920";
    tmp(42786) := x"0920";
    tmp(42787) := x"0920";
    tmp(42788) := x"0920";
    tmp(42789) := x"0920";
    tmp(42790) := x"0920";
    tmp(42791) := x"0920";
    tmp(42792) := x"0920";
    tmp(42793) := x"0920";
    tmp(42794) := x"0900";
    tmp(42795) := x"0900";
    tmp(42796) := x"0900";
    tmp(42797) := x"0900";
    tmp(42798) := x"0900";
    tmp(42799) := x"0900";
    tmp(42800) := x"0900";
    tmp(42801) := x"0900";
    tmp(42802) := x"0900";
    tmp(42803) := x"0900";
    tmp(42804) := x"0900";
    tmp(42805) := x"0900";
    tmp(42806) := x"0900";
    tmp(42807) := x"0900";
    tmp(42808) := x"0900";
    tmp(42809) := x"0900";
    tmp(42810) := x"0900";
    tmp(42811) := x"0900";
    tmp(42812) := x"0900";
    tmp(42813) := x"0900";
    tmp(42814) := x"0920";
    tmp(42815) := x"0920";
    tmp(42816) := x"0920";
    tmp(42817) := x"0920";
    tmp(42818) := x"0920";
    tmp(42819) := x"0920";
    tmp(42820) := x"0920";
    tmp(42821) := x"0920";
    tmp(42822) := x"0900";
    tmp(42823) := x"0900";
    tmp(42824) := x"0900";
    tmp(42825) := x"08e0";
    tmp(42826) := x"08e0";
    tmp(42827) := x"08e0";
    tmp(42828) := x"08e0";
    tmp(42829) := x"08c0";
    tmp(42830) := x"08c0";
    tmp(42831) := x"08a0";
    tmp(42832) := x"08a0";
    tmp(42833) := x"2101";
    tmp(42834) := x"6203";
    tmp(42835) := x"8a65";
    tmp(42836) := x"9a86";
    tmp(42837) := x"9aa7";
    tmp(42838) := x"aae9";
    tmp(42839) := x"b2e9";
    tmp(42840) := x"bb2a";
    tmp(42841) := x"c36b";
    tmp(42842) := x"cb8c";
    tmp(42843) := x"cb6c";
    tmp(42844) := x"cb6b";
    tmp(42845) := x"d36b";
    tmp(42846) := x"c309";
    tmp(42847) := x"cb09";
    tmp(42848) := x"cb09";
    tmp(42849) := x"c2e9";
    tmp(42850) := x"b2c8";
    tmp(42851) := x"dc0d";
    tmp(42852) := x"cb8c";
    tmp(42853) := x"d38b";
    tmp(42854) := x"dbab";
    tmp(42855) := x"cb6a";
    tmp(42856) := x"dbab";
    tmp(42857) := x"e3cb";
    tmp(42858) := x"e3cb";
    tmp(42859) := x"e3cc";
    tmp(42860) := x"dbcc";
    tmp(42861) := x"f48e";
    tmp(42862) := x"f531";
    tmp(42863) := x"fcf1";
    tmp(42864) := x"fccf";
    tmp(42865) := x"fcf0";
    tmp(42866) := x"f4b0";
    tmp(42867) := x"fcd1";
    tmp(42868) := x"fd12";
    tmp(42869) := x"fcf2";
    tmp(42870) := x"f4d2";
    tmp(42871) := x"ec72";
    tmp(42872) := x"e471";
    tmp(42873) := x"ec72";
    tmp(42874) := x"d3ae";
    tmp(42875) := x"9206";
    tmp(42876) := x"4061";
    tmp(42877) := x"2020";
    tmp(42878) := x"1000";
    tmp(42879) := x"0800";
    tmp(42880) := x"0800";
    tmp(42881) := x"1000";
    tmp(42882) := x"0800";
    tmp(42883) := x"1000";
    tmp(42884) := x"1800";
    tmp(42885) := x"3000";
    tmp(42886) := x"3800";
    tmp(42887) := x"3000";
    tmp(42888) := x"3000";
    tmp(42889) := x"4000";
    tmp(42890) := x"5000";
    tmp(42891) := x"7000";
    tmp(42892) := x"8820";
    tmp(42893) := x"9020";
    tmp(42894) := x"a821";
    tmp(42895) := x"c041";
    tmp(42896) := x"e061";
    tmp(42897) := x"5861";
    tmp(42898) := x"1040";
    tmp(42899) := x"1040";
    tmp(42900) := x"1040";
    tmp(42901) := x"0840";
    tmp(42902) := x"0840";
    tmp(42903) := x"0840";
    tmp(42904) := x"0840";
    tmp(42905) := x"0840";
    tmp(42906) := x"0840";
    tmp(42907) := x"0840";
    tmp(42908) := x"0840";
    tmp(42909) := x"0840";
    tmp(42910) := x"0840";
    tmp(42911) := x"0840";
    tmp(42912) := x"0840";
    tmp(42913) := x"0840";
    tmp(42914) := x"0840";
    tmp(42915) := x"0840";
    tmp(42916) := x"0840";
    tmp(42917) := x"001f";
    tmp(42918) := x"001f";
    tmp(42919) := x"001f";
    tmp(42920) := x"001f";
    tmp(42921) := x"001f";
    tmp(42922) := x"001f";
    tmp(42923) := x"001f";
    tmp(42924) := x"001f";
    tmp(42925) := x"001f";
    tmp(42926) := x"001f";
    tmp(42927) := x"001f";
    tmp(42928) := x"001f";
    tmp(42929) := x"001f";
    tmp(42930) := x"001f";
    tmp(42931) := x"001f";
    tmp(42932) := x"001f";
    tmp(42933) := x"001f";
    tmp(42934) := x"001f";
    tmp(42935) := x"001f";
    tmp(42936) := x"001f";
    tmp(42937) := x"001f";
    tmp(42938) := x"001f";
    tmp(42939) := x"001f";
    tmp(42940) := x"001f";
    tmp(42941) := x"001f";
    tmp(42942) := x"001f";
    tmp(42943) := x"001f";
    tmp(42944) := x"001f";
    tmp(42945) := x"001f";
    tmp(42946) := x"001f";
    tmp(42947) := x"001f";
    tmp(42948) := x"001f";
    tmp(42949) := x"001f";
    tmp(42950) := x"001f";
    tmp(42951) := x"001f";
    tmp(42952) := x"001f";
    tmp(42953) := x"001f";
    tmp(42954) := x"001f";
    tmp(42955) := x"001f";
    tmp(42956) := x"001f";
    tmp(42957) := x"1061";
    tmp(42958) := x"1061";
    tmp(42959) := x"1061";
    tmp(42960) := x"0000";
    tmp(42961) := x"0880";
    tmp(42962) := x"0880";
    tmp(42963) := x"0880";
    tmp(42964) := x"0880";
    tmp(42965) := x"0880";
    tmp(42966) := x"0880";
    tmp(42967) := x"0860";
    tmp(42968) := x"0860";
    tmp(42969) := x"0860";
    tmp(42970) := x"0860";
    tmp(42971) := x"0860";
    tmp(42972) := x"0840";
    tmp(42973) := x"0840";
    tmp(42974) := x"0840";
    tmp(42975) := x"0840";
    tmp(42976) := x"0840";
    tmp(42977) := x"0840";
    tmp(42978) := x"0840";
    tmp(42979) := x"0840";
    tmp(42980) := x"0840";
    tmp(42981) := x"0840";
    tmp(42982) := x"0840";
    tmp(42983) := x"0840";
    tmp(42984) := x"0860";
    tmp(42985) := x"0860";
    tmp(42986) := x"0860";
    tmp(42987) := x"0860";
    tmp(42988) := x"0880";
    tmp(42989) := x"08a0";
    tmp(42990) := x"08a0";
    tmp(42991) := x"08a0";
    tmp(42992) := x"08a0";
    tmp(42993) := x"08a0";
    tmp(42994) := x"08c0";
    tmp(42995) := x"08c0";
    tmp(42996) := x"08c0";
    tmp(42997) := x"08c0";
    tmp(42998) := x"08c0";
    tmp(42999) := x"08e0";
    tmp(43000) := x"08e0";
    tmp(43001) := x"0900";
    tmp(43002) := x"0900";
    tmp(43003) := x"0900";
    tmp(43004) := x"0900";
    tmp(43005) := x"0900";
    tmp(43006) := x"0900";
    tmp(43007) := x"0900";
    tmp(43008) := x"0900";
    tmp(43009) := x"0900";
    tmp(43010) := x"0900";
    tmp(43011) := x"0900";
    tmp(43012) := x"0920";
    tmp(43013) := x"0920";
    tmp(43014) := x"0920";
    tmp(43015) := x"0920";
    tmp(43016) := x"0920";
    tmp(43017) := x"0920";
    tmp(43018) := x"0940";
    tmp(43019) := x"0920";
    tmp(43020) := x"0920";
    tmp(43021) := x"0920";
    tmp(43022) := x"0920";
    tmp(43023) := x"0920";
    tmp(43024) := x"0920";
    tmp(43025) := x"0920";
    tmp(43026) := x"0920";
    tmp(43027) := x"0900";
    tmp(43028) := x"0920";
    tmp(43029) := x"0920";
    tmp(43030) := x"0920";
    tmp(43031) := x"0920";
    tmp(43032) := x"0920";
    tmp(43033) := x"0920";
    tmp(43034) := x"0900";
    tmp(43035) := x"0900";
    tmp(43036) := x"0900";
    tmp(43037) := x"0900";
    tmp(43038) := x"0900";
    tmp(43039) := x"0900";
    tmp(43040) := x"0900";
    tmp(43041) := x"0900";
    tmp(43042) := x"0900";
    tmp(43043) := x"0900";
    tmp(43044) := x"0900";
    tmp(43045) := x"0900";
    tmp(43046) := x"0900";
    tmp(43047) := x"0900";
    tmp(43048) := x"0900";
    tmp(43049) := x"0900";
    tmp(43050) := x"0900";
    tmp(43051) := x"0900";
    tmp(43052) := x"0900";
    tmp(43053) := x"0920";
    tmp(43054) := x"0920";
    tmp(43055) := x"0920";
    tmp(43056) := x"0920";
    tmp(43057) := x"0920";
    tmp(43058) := x"0920";
    tmp(43059) := x"0920";
    tmp(43060) := x"0920";
    tmp(43061) := x"0920";
    tmp(43062) := x"0900";
    tmp(43063) := x"0900";
    tmp(43064) := x"0900";
    tmp(43065) := x"08e0";
    tmp(43066) := x"08e0";
    tmp(43067) := x"08e0";
    tmp(43068) := x"08c0";
    tmp(43069) := x"08c0";
    tmp(43070) := x"08a0";
    tmp(43071) := x"10c0";
    tmp(43072) := x"3161";
    tmp(43073) := x"7244";
    tmp(43074) := x"8a44";
    tmp(43075) := x"9266";
    tmp(43076) := x"aae8";
    tmp(43077) := x"b34a";
    tmp(43078) := x"b34b";
    tmp(43079) := x"bb4b";
    tmp(43080) := x"cb8c";
    tmp(43081) := x"c38b";
    tmp(43082) := x"cb8c";
    tmp(43083) := x"d3ad";
    tmp(43084) := x"cb8c";
    tmp(43085) := x"db8b";
    tmp(43086) := x"d34a";
    tmp(43087) := x"cb2a";
    tmp(43088) := x"c2c9";
    tmp(43089) := x"bac9";
    tmp(43090) := x"cb4a";
    tmp(43091) := x"d38b";
    tmp(43092) := x"bb2a";
    tmp(43093) := x"cb6b";
    tmp(43094) := x"cb4a";
    tmp(43095) := x"c349";
    tmp(43096) := x"dbab";
    tmp(43097) := x"dbab";
    tmp(43098) := x"dbcb";
    tmp(43099) := x"dbcc";
    tmp(43100) := x"ec2e";
    tmp(43101) := x"e40e";
    tmp(43102) := x"dbee";
    tmp(43103) := x"e42e";
    tmp(43104) := x"ec4d";
    tmp(43105) := x"fcaf";
    tmp(43106) := x"ec6f";
    tmp(43107) := x"f4d0";
    tmp(43108) := x"f4d1";
    tmp(43109) := x"f4d1";
    tmp(43110) := x"f4d2";
    tmp(43111) := x"ec51";
    tmp(43112) := x"e452";
    tmp(43113) := x"dc31";
    tmp(43114) := x"bb2c";
    tmp(43115) := x"89e6";
    tmp(43116) := x"60e3";
    tmp(43117) := x"3841";
    tmp(43118) := x"1000";
    tmp(43119) := x"0800";
    tmp(43120) := x"0800";
    tmp(43121) := x"0800";
    tmp(43122) := x"0800";
    tmp(43123) := x"1000";
    tmp(43124) := x"1800";
    tmp(43125) := x"3000";
    tmp(43126) := x"3800";
    tmp(43127) := x"3000";
    tmp(43128) := x"3800";
    tmp(43129) := x"5000";
    tmp(43130) := x"5800";
    tmp(43131) := x"6800";
    tmp(43132) := x"8020";
    tmp(43133) := x"9020";
    tmp(43134) := x"a841";
    tmp(43135) := x"d861";
    tmp(43136) := x"c841";
    tmp(43137) := x"c061";
    tmp(43138) := x"3041";
    tmp(43139) := x"1040";
    tmp(43140) := x"1040";
    tmp(43141) := x"0840";
    tmp(43142) := x"0840";
    tmp(43143) := x"0840";
    tmp(43144) := x"0840";
    tmp(43145) := x"0840";
    tmp(43146) := x"0840";
    tmp(43147) := x"0840";
    tmp(43148) := x"0840";
    tmp(43149) := x"0840";
    tmp(43150) := x"0840";
    tmp(43151) := x"0840";
    tmp(43152) := x"0840";
    tmp(43153) := x"0840";
    tmp(43154) := x"0840";
    tmp(43155) := x"0840";
    tmp(43156) := x"0840";
    tmp(43157) := x"001f";
    tmp(43158) := x"001f";
    tmp(43159) := x"001f";
    tmp(43160) := x"001f";
    tmp(43161) := x"001f";
    tmp(43162) := x"001f";
    tmp(43163) := x"001f";
    tmp(43164) := x"001f";
    tmp(43165) := x"001f";
    tmp(43166) := x"001f";
    tmp(43167) := x"001f";
    tmp(43168) := x"001f";
    tmp(43169) := x"001f";
    tmp(43170) := x"001f";
    tmp(43171) := x"001f";
    tmp(43172) := x"001f";
    tmp(43173) := x"001f";
    tmp(43174) := x"001f";
    tmp(43175) := x"001f";
    tmp(43176) := x"001f";
    tmp(43177) := x"001f";
    tmp(43178) := x"001f";
    tmp(43179) := x"001f";
    tmp(43180) := x"001f";
    tmp(43181) := x"001f";
    tmp(43182) := x"001f";
    tmp(43183) := x"001f";
    tmp(43184) := x"001f";
    tmp(43185) := x"001f";
    tmp(43186) := x"001f";
    tmp(43187) := x"001f";
    tmp(43188) := x"001f";
    tmp(43189) := x"001f";
    tmp(43190) := x"001f";
    tmp(43191) := x"001f";
    tmp(43192) := x"001f";
    tmp(43193) := x"001f";
    tmp(43194) := x"001f";
    tmp(43195) := x"001f";
    tmp(43196) := x"001f";
    tmp(43197) := x"1061";
    tmp(43198) := x"1061";
    tmp(43199) := x"1061";
    tmp(43200) := x"0000";
    tmp(43201) := x"08a0";
    tmp(43202) := x"0880";
    tmp(43203) := x"0880";
    tmp(43204) := x"0880";
    tmp(43205) := x"0880";
    tmp(43206) := x"0880";
    tmp(43207) := x"0860";
    tmp(43208) := x"0860";
    tmp(43209) := x"0860";
    tmp(43210) := x"0860";
    tmp(43211) := x"0860";
    tmp(43212) := x"0860";
    tmp(43213) := x"0840";
    tmp(43214) := x"0840";
    tmp(43215) := x"0840";
    tmp(43216) := x"0840";
    tmp(43217) := x"0840";
    tmp(43218) := x"0840";
    tmp(43219) := x"0840";
    tmp(43220) := x"0840";
    tmp(43221) := x"0840";
    tmp(43222) := x"0840";
    tmp(43223) := x"0840";
    tmp(43224) := x"0840";
    tmp(43225) := x"0840";
    tmp(43226) := x"0860";
    tmp(43227) := x"0860";
    tmp(43228) := x"0860";
    tmp(43229) := x"0880";
    tmp(43230) := x"08a0";
    tmp(43231) := x"08a0";
    tmp(43232) := x"08a0";
    tmp(43233) := x"08a0";
    tmp(43234) := x"08a0";
    tmp(43235) := x"08c0";
    tmp(43236) := x"08c0";
    tmp(43237) := x"08c0";
    tmp(43238) := x"08c0";
    tmp(43239) := x"08e0";
    tmp(43240) := x"08e0";
    tmp(43241) := x"0900";
    tmp(43242) := x"0900";
    tmp(43243) := x"0900";
    tmp(43244) := x"0900";
    tmp(43245) := x"0900";
    tmp(43246) := x"0900";
    tmp(43247) := x"0900";
    tmp(43248) := x"0900";
    tmp(43249) := x"0900";
    tmp(43250) := x"0900";
    tmp(43251) := x"0900";
    tmp(43252) := x"0900";
    tmp(43253) := x"0920";
    tmp(43254) := x"0920";
    tmp(43255) := x"0920";
    tmp(43256) := x"0920";
    tmp(43257) := x"0920";
    tmp(43258) := x"0920";
    tmp(43259) := x"0920";
    tmp(43260) := x"0920";
    tmp(43261) := x"0920";
    tmp(43262) := x"0920";
    tmp(43263) := x"0920";
    tmp(43264) := x"0920";
    tmp(43265) := x"0920";
    tmp(43266) := x"0920";
    tmp(43267) := x"0900";
    tmp(43268) := x"0900";
    tmp(43269) := x"0900";
    tmp(43270) := x"0900";
    tmp(43271) := x"0920";
    tmp(43272) := x"0900";
    tmp(43273) := x"0900";
    tmp(43274) := x"0900";
    tmp(43275) := x"0900";
    tmp(43276) := x"0900";
    tmp(43277) := x"0900";
    tmp(43278) := x"0900";
    tmp(43279) := x"0900";
    tmp(43280) := x"0900";
    tmp(43281) := x"0900";
    tmp(43282) := x"0900";
    tmp(43283) := x"0900";
    tmp(43284) := x"0900";
    tmp(43285) := x"0900";
    tmp(43286) := x"0900";
    tmp(43287) := x"0900";
    tmp(43288) := x"0900";
    tmp(43289) := x"0900";
    tmp(43290) := x"0900";
    tmp(43291) := x"0900";
    tmp(43292) := x"0900";
    tmp(43293) := x"0900";
    tmp(43294) := x"0920";
    tmp(43295) := x"0920";
    tmp(43296) := x"0920";
    tmp(43297) := x"0920";
    tmp(43298) := x"0920";
    tmp(43299) := x"0920";
    tmp(43300) := x"0920";
    tmp(43301) := x"0920";
    tmp(43302) := x"0900";
    tmp(43303) := x"0900";
    tmp(43304) := x"0900";
    tmp(43305) := x"0900";
    tmp(43306) := x"08e0";
    tmp(43307) := x"08e0";
    tmp(43308) := x"08c0";
    tmp(43309) := x"08a0";
    tmp(43310) := x"18e0";
    tmp(43311) := x"4181";
    tmp(43312) := x"8244";
    tmp(43313) := x"8224";
    tmp(43314) := x"8a25";
    tmp(43315) := x"a2c8";
    tmp(43316) := x"bb4b";
    tmp(43317) := x"c38d";
    tmp(43318) := x"c3ad";
    tmp(43319) := x"cbad";
    tmp(43320) := x"c3ad";
    tmp(43321) := x"c3ad";
    tmp(43322) := x"cb8c";
    tmp(43323) := x"cb6c";
    tmp(43324) := x"cb6c";
    tmp(43325) := x"cb4b";
    tmp(43326) := x"cb4a";
    tmp(43327) := x"c2ea";
    tmp(43328) := x"baa9";
    tmp(43329) := x"b2c9";
    tmp(43330) := x"d38c";
    tmp(43331) := x"cb4b";
    tmp(43332) := x"c34a";
    tmp(43333) := x"d38c";
    tmp(43334) := x"cb4b";
    tmp(43335) := x"c34a";
    tmp(43336) := x"d38b";
    tmp(43337) := x"dbcc";
    tmp(43338) := x"dbab";
    tmp(43339) := x"dbec";
    tmp(43340) := x"e3ed";
    tmp(43341) := x"d38c";
    tmp(43342) := x"e40e";
    tmp(43343) := x"ec6f";
    tmp(43344) := x"dc0d";
    tmp(43345) := x"f490";
    tmp(43346) := x"ec90";
    tmp(43347) := x"ecb0";
    tmp(43348) := x"e46f";
    tmp(43349) := x"ecb1";
    tmp(43350) := x"dc4f";
    tmp(43351) := x"e491";
    tmp(43352) := x"dc52";
    tmp(43353) := x"cbf0";
    tmp(43354) := x"a2aa";
    tmp(43355) := x"7965";
    tmp(43356) := x"7124";
    tmp(43357) := x"58e3";
    tmp(43358) := x"2020";
    tmp(43359) := x"0800";
    tmp(43360) := x"0800";
    tmp(43361) := x"0800";
    tmp(43362) := x"0800";
    tmp(43363) := x"1000";
    tmp(43364) := x"1800";
    tmp(43365) := x"2800";
    tmp(43366) := x"3800";
    tmp(43367) := x"4000";
    tmp(43368) := x"4800";
    tmp(43369) := x"5000";
    tmp(43370) := x"5000";
    tmp(43371) := x"6000";
    tmp(43372) := x"8020";
    tmp(43373) := x"8820";
    tmp(43374) := x"9020";
    tmp(43375) := x"b841";
    tmp(43376) := x"e061";
    tmp(43377) := x"c841";
    tmp(43378) := x"a081";
    tmp(43379) := x"2040";
    tmp(43380) := x"1040";
    tmp(43381) := x"1040";
    tmp(43382) := x"0840";
    tmp(43383) := x"0840";
    tmp(43384) := x"0840";
    tmp(43385) := x"0840";
    tmp(43386) := x"0840";
    tmp(43387) := x"0840";
    tmp(43388) := x"0840";
    tmp(43389) := x"0840";
    tmp(43390) := x"0840";
    tmp(43391) := x"0840";
    tmp(43392) := x"0840";
    tmp(43393) := x"0840";
    tmp(43394) := x"0840";
    tmp(43395) := x"0840";
    tmp(43396) := x"0840";
    tmp(43397) := x"001f";
    tmp(43398) := x"001f";
    tmp(43399) := x"001f";
    tmp(43400) := x"001f";
    tmp(43401) := x"001f";
    tmp(43402) := x"001f";
    tmp(43403) := x"001f";
    tmp(43404) := x"001f";
    tmp(43405) := x"001f";
    tmp(43406) := x"001f";
    tmp(43407) := x"001f";
    tmp(43408) := x"001f";
    tmp(43409) := x"001f";
    tmp(43410) := x"001f";
    tmp(43411) := x"001f";
    tmp(43412) := x"001f";
    tmp(43413) := x"001f";
    tmp(43414) := x"001f";
    tmp(43415) := x"001f";
    tmp(43416) := x"001f";
    tmp(43417) := x"001f";
    tmp(43418) := x"001f";
    tmp(43419) := x"001f";
    tmp(43420) := x"001f";
    tmp(43421) := x"001f";
    tmp(43422) := x"001f";
    tmp(43423) := x"001f";
    tmp(43424) := x"001f";
    tmp(43425) := x"001f";
    tmp(43426) := x"001f";
    tmp(43427) := x"001f";
    tmp(43428) := x"001f";
    tmp(43429) := x"001f";
    tmp(43430) := x"001f";
    tmp(43431) := x"001f";
    tmp(43432) := x"001f";
    tmp(43433) := x"001f";
    tmp(43434) := x"001f";
    tmp(43435) := x"001f";
    tmp(43436) := x"001f";
    tmp(43437) := x"1060";
    tmp(43438) := x"1061";
    tmp(43439) := x"1061";
    tmp(43440) := x"0000";
    tmp(43441) := x"08a0";
    tmp(43442) := x"0880";
    tmp(43443) := x"0880";
    tmp(43444) := x"0880";
    tmp(43445) := x"0880";
    tmp(43446) := x"0880";
    tmp(43447) := x"0880";
    tmp(43448) := x"0860";
    tmp(43449) := x"0860";
    tmp(43450) := x"0860";
    tmp(43451) := x"0860";
    tmp(43452) := x"0860";
    tmp(43453) := x"0860";
    tmp(43454) := x"0840";
    tmp(43455) := x"0840";
    tmp(43456) := x"0840";
    tmp(43457) := x"0840";
    tmp(43458) := x"0840";
    tmp(43459) := x"0840";
    tmp(43460) := x"0840";
    tmp(43461) := x"0840";
    tmp(43462) := x"0840";
    tmp(43463) := x"0840";
    tmp(43464) := x"0840";
    tmp(43465) := x"0840";
    tmp(43466) := x"0840";
    tmp(43467) := x"0860";
    tmp(43468) := x"0860";
    tmp(43469) := x"0860";
    tmp(43470) := x"0880";
    tmp(43471) := x"08a0";
    tmp(43472) := x"08a0";
    tmp(43473) := x"08a0";
    tmp(43474) := x"08a0";
    tmp(43475) := x"08a0";
    tmp(43476) := x"08a0";
    tmp(43477) := x"08c0";
    tmp(43478) := x"08c0";
    tmp(43479) := x"08c0";
    tmp(43480) := x"08c0";
    tmp(43481) := x"08e0";
    tmp(43482) := x"0900";
    tmp(43483) := x"08e0";
    tmp(43484) := x"0900";
    tmp(43485) := x"0900";
    tmp(43486) := x"0900";
    tmp(43487) := x"0900";
    tmp(43488) := x"0900";
    tmp(43489) := x"0900";
    tmp(43490) := x"0900";
    tmp(43491) := x"0900";
    tmp(43492) := x"0900";
    tmp(43493) := x"0900";
    tmp(43494) := x"0920";
    tmp(43495) := x"0920";
    tmp(43496) := x"0920";
    tmp(43497) := x"0920";
    tmp(43498) := x"0920";
    tmp(43499) := x"0920";
    tmp(43500) := x"0920";
    tmp(43501) := x"0920";
    tmp(43502) := x"0920";
    tmp(43503) := x"0920";
    tmp(43504) := x"0920";
    tmp(43505) := x"0920";
    tmp(43506) := x"0900";
    tmp(43507) := x"0900";
    tmp(43508) := x"0900";
    tmp(43509) := x"0900";
    tmp(43510) := x"0900";
    tmp(43511) := x"0900";
    tmp(43512) := x"0900";
    tmp(43513) := x"0900";
    tmp(43514) := x"0900";
    tmp(43515) := x"0900";
    tmp(43516) := x"0900";
    tmp(43517) := x"08e0";
    tmp(43518) := x"0900";
    tmp(43519) := x"08e0";
    tmp(43520) := x"08e0";
    tmp(43521) := x"0900";
    tmp(43522) := x"0900";
    tmp(43523) := x"08e0";
    tmp(43524) := x"08e0";
    tmp(43525) := x"0900";
    tmp(43526) := x"0900";
    tmp(43527) := x"0900";
    tmp(43528) := x"0900";
    tmp(43529) := x"0900";
    tmp(43530) := x"0900";
    tmp(43531) := x"0900";
    tmp(43532) := x"0900";
    tmp(43533) := x"0920";
    tmp(43534) := x"0920";
    tmp(43535) := x"0920";
    tmp(43536) := x"0920";
    tmp(43537) := x"0920";
    tmp(43538) := x"0920";
    tmp(43539) := x"0920";
    tmp(43540) := x"0920";
    tmp(43541) := x"0920";
    tmp(43542) := x"0920";
    tmp(43543) := x"0900";
    tmp(43544) := x"0900";
    tmp(43545) := x"08e0";
    tmp(43546) := x"08e0";
    tmp(43547) := x"08e0";
    tmp(43548) := x"08a0";
    tmp(43549) := x"1900";
    tmp(43550) := x"51a2";
    tmp(43551) := x"7a04";
    tmp(43552) := x"8a25";
    tmp(43553) := x"9246";
    tmp(43554) := x"a2c8";
    tmp(43555) := x"ab4b";
    tmp(43556) := x"c3cf";
    tmp(43557) := x"cbef";
    tmp(43558) := x"d42f";
    tmp(43559) := x"dc0f";
    tmp(43560) := x"cbce";
    tmp(43561) := x"cbae";
    tmp(43562) := x"c36d";
    tmp(43563) := x"cb6c";
    tmp(43564) := x"cb6c";
    tmp(43565) := x"cb6c";
    tmp(43566) := x"c32a";
    tmp(43567) := x"c2c9";
    tmp(43568) := x"b2a9";
    tmp(43569) := x"c34b";
    tmp(43570) := x"d3ad";
    tmp(43571) := x"c34b";
    tmp(43572) := x"cb2b";
    tmp(43573) := x"d3ac";
    tmp(43574) := x"d38b";
    tmp(43575) := x"c329";
    tmp(43576) := x"cb4a";
    tmp(43577) := x"d36a";
    tmp(43578) := x"db8a";
    tmp(43579) := x"dbec";
    tmp(43580) := x"dbed";
    tmp(43581) := x"d3cc";
    tmp(43582) := x"e44e";
    tmp(43583) := x"ec4e";
    tmp(43584) := x"d3ed";
    tmp(43585) := x"d40e";
    tmp(43586) := x"d40e";
    tmp(43587) := x"bb8d";
    tmp(43588) := x"bb4c";
    tmp(43589) := x"bb8d";
    tmp(43590) := x"bb6d";
    tmp(43591) := x"c3ef";
    tmp(43592) := x"c3cf";
    tmp(43593) := x"b34d";
    tmp(43594) := x"8a28";
    tmp(43595) := x"7104";
    tmp(43596) := x"58c3";
    tmp(43597) := x"58e3";
    tmp(43598) := x"2841";
    tmp(43599) := x"0800";
    tmp(43600) := x"0800";
    tmp(43601) := x"0800";
    tmp(43602) := x"0800";
    tmp(43603) := x"1000";
    tmp(43604) := x"1800";
    tmp(43605) := x"2800";
    tmp(43606) := x"3800";
    tmp(43607) := x"4800";
    tmp(43608) := x"5000";
    tmp(43609) := x"5000";
    tmp(43610) := x"5000";
    tmp(43611) := x"5800";
    tmp(43612) := x"6800";
    tmp(43613) := x"7820";
    tmp(43614) := x"8020";
    tmp(43615) := x"8020";
    tmp(43616) := x"b021";
    tmp(43617) := x"d041";
    tmp(43618) := x"f061";
    tmp(43619) := x"8881";
    tmp(43620) := x"2040";
    tmp(43621) := x"1040";
    tmp(43622) := x"0840";
    tmp(43623) := x"0840";
    tmp(43624) := x"0840";
    tmp(43625) := x"0840";
    tmp(43626) := x"0840";
    tmp(43627) := x"0840";
    tmp(43628) := x"0840";
    tmp(43629) := x"0840";
    tmp(43630) := x"0840";
    tmp(43631) := x"0840";
    tmp(43632) := x"0840";
    tmp(43633) := x"0840";
    tmp(43634) := x"0840";
    tmp(43635) := x"0840";
    tmp(43636) := x"0840";
    tmp(43637) := x"001f";
    tmp(43638) := x"001f";
    tmp(43639) := x"001f";
    tmp(43640) := x"001f";
    tmp(43641) := x"001f";
    tmp(43642) := x"001f";
    tmp(43643) := x"001f";
    tmp(43644) := x"001f";
    tmp(43645) := x"001f";
    tmp(43646) := x"001f";
    tmp(43647) := x"001f";
    tmp(43648) := x"001f";
    tmp(43649) := x"001f";
    tmp(43650) := x"001f";
    tmp(43651) := x"001f";
    tmp(43652) := x"001f";
    tmp(43653) := x"001f";
    tmp(43654) := x"001f";
    tmp(43655) := x"001f";
    tmp(43656) := x"001f";
    tmp(43657) := x"001f";
    tmp(43658) := x"001f";
    tmp(43659) := x"001f";
    tmp(43660) := x"001f";
    tmp(43661) := x"001f";
    tmp(43662) := x"001f";
    tmp(43663) := x"001f";
    tmp(43664) := x"001f";
    tmp(43665) := x"001f";
    tmp(43666) := x"001f";
    tmp(43667) := x"001f";
    tmp(43668) := x"001f";
    tmp(43669) := x"001f";
    tmp(43670) := x"001f";
    tmp(43671) := x"001f";
    tmp(43672) := x"001f";
    tmp(43673) := x"001f";
    tmp(43674) := x"001f";
    tmp(43675) := x"001f";
    tmp(43676) := x"001f";
    tmp(43677) := x"1060";
    tmp(43678) := x"1061";
    tmp(43679) := x"1061";
    tmp(43680) := x"0000";
    tmp(43681) := x"0880";
    tmp(43682) := x"0880";
    tmp(43683) := x"0880";
    tmp(43684) := x"0880";
    tmp(43685) := x"0880";
    tmp(43686) := x"0880";
    tmp(43687) := x"0880";
    tmp(43688) := x"0880";
    tmp(43689) := x"0860";
    tmp(43690) := x"0860";
    tmp(43691) := x"0860";
    tmp(43692) := x"0860";
    tmp(43693) := x"0860";
    tmp(43694) := x"0860";
    tmp(43695) := x"0860";
    tmp(43696) := x"0840";
    tmp(43697) := x"0840";
    tmp(43698) := x"0840";
    tmp(43699) := x"0840";
    tmp(43700) := x"0840";
    tmp(43701) := x"0840";
    tmp(43702) := x"0840";
    tmp(43703) := x"0840";
    tmp(43704) := x"0840";
    tmp(43705) := x"0840";
    tmp(43706) := x"0840";
    tmp(43707) := x"0840";
    tmp(43708) := x"0840";
    tmp(43709) := x"0860";
    tmp(43710) := x"0860";
    tmp(43711) := x"0880";
    tmp(43712) := x"0880";
    tmp(43713) := x"08a0";
    tmp(43714) := x"08a0";
    tmp(43715) := x"08a0";
    tmp(43716) := x"08a0";
    tmp(43717) := x"08a0";
    tmp(43718) := x"08a0";
    tmp(43719) := x"08c0";
    tmp(43720) := x"08c0";
    tmp(43721) := x"08e0";
    tmp(43722) := x"08e0";
    tmp(43723) := x"08e0";
    tmp(43724) := x"0900";
    tmp(43725) := x"0900";
    tmp(43726) := x"08e0";
    tmp(43727) := x"0900";
    tmp(43728) := x"0900";
    tmp(43729) := x"0900";
    tmp(43730) := x"0900";
    tmp(43731) := x"0900";
    tmp(43732) := x"0900";
    tmp(43733) := x"0900";
    tmp(43734) := x"0900";
    tmp(43735) := x"0920";
    tmp(43736) := x"0920";
    tmp(43737) := x"0920";
    tmp(43738) := x"0920";
    tmp(43739) := x"0920";
    tmp(43740) := x"0920";
    tmp(43741) := x"0920";
    tmp(43742) := x"0920";
    tmp(43743) := x"0920";
    tmp(43744) := x"0920";
    tmp(43745) := x"0920";
    tmp(43746) := x"0900";
    tmp(43747) := x"0900";
    tmp(43748) := x"0900";
    tmp(43749) := x"0900";
    tmp(43750) := x"0900";
    tmp(43751) := x"0900";
    tmp(43752) := x"0900";
    tmp(43753) := x"0900";
    tmp(43754) := x"0900";
    tmp(43755) := x"0900";
    tmp(43756) := x"0900";
    tmp(43757) := x"08e0";
    tmp(43758) := x"0900";
    tmp(43759) := x"08e0";
    tmp(43760) := x"08e0";
    tmp(43761) := x"08e0";
    tmp(43762) := x"08e0";
    tmp(43763) := x"08e0";
    tmp(43764) := x"08e0";
    tmp(43765) := x"0900";
    tmp(43766) := x"0900";
    tmp(43767) := x"0900";
    tmp(43768) := x"0900";
    tmp(43769) := x"0900";
    tmp(43770) := x"0900";
    tmp(43771) := x"0900";
    tmp(43772) := x"0920";
    tmp(43773) := x"0920";
    tmp(43774) := x"0920";
    tmp(43775) := x"0920";
    tmp(43776) := x"0920";
    tmp(43777) := x"0920";
    tmp(43778) := x"0920";
    tmp(43779) := x"0920";
    tmp(43780) := x"0920";
    tmp(43781) := x"0920";
    tmp(43782) := x"0900";
    tmp(43783) := x"0900";
    tmp(43784) := x"0900";
    tmp(43785) := x"08e0";
    tmp(43786) := x"08e0";
    tmp(43787) := x"08c0";
    tmp(43788) := x"1900";
    tmp(43789) := x"51a2";
    tmp(43790) := x"79e3";
    tmp(43791) := x"8224";
    tmp(43792) := x"8a46";
    tmp(43793) := x"9aa9";
    tmp(43794) := x"b34c";
    tmp(43795) := x"c3cf";
    tmp(43796) := x"cc71";
    tmp(43797) := x"d451";
    tmp(43798) := x"dc71";
    tmp(43799) := x"d430";
    tmp(43800) := x"c3ae";
    tmp(43801) := x"cbae";
    tmp(43802) := x"c36c";
    tmp(43803) := x"cbcd";
    tmp(43804) := x"cb8d";
    tmp(43805) := x"cb6c";
    tmp(43806) := x"baea";
    tmp(43807) := x"b289";
    tmp(43808) := x"baea";
    tmp(43809) := x"cbad";
    tmp(43810) := x"cb8c";
    tmp(43811) := x"bb0a";
    tmp(43812) := x"cb4b";
    tmp(43813) := x"cb6b";
    tmp(43814) := x"c32a";
    tmp(43815) := x"c329";
    tmp(43816) := x"cb49";
    tmp(43817) := x"cb49";
    tmp(43818) := x"d38a";
    tmp(43819) := x"cb6a";
    tmp(43820) := x"cb6a";
    tmp(43821) := x"c36a";
    tmp(43822) := x"aae9";
    tmp(43823) := x"b309";
    tmp(43824) := x"9aa9";
    tmp(43825) := x"9ac9";
    tmp(43826) := x"8a68";
    tmp(43827) := x"8a48";
    tmp(43828) := x"8227";
    tmp(43829) := x"71e7";
    tmp(43830) := x"69c7";
    tmp(43831) := x"5986";
    tmp(43832) := x"59a6";
    tmp(43833) := x"5166";
    tmp(43834) := x"5924";
    tmp(43835) := x"8165";
    tmp(43836) := x"6904";
    tmp(43837) := x"50c3";
    tmp(43838) := x"2021";
    tmp(43839) := x"0800";
    tmp(43840) := x"1000";
    tmp(43841) := x"1000";
    tmp(43842) := x"0800";
    tmp(43843) := x"1000";
    tmp(43844) := x"1800";
    tmp(43845) := x"2000";
    tmp(43846) := x"3800";
    tmp(43847) := x"4800";
    tmp(43848) := x"5000";
    tmp(43849) := x"5800";
    tmp(43850) := x"5800";
    tmp(43851) := x"5800";
    tmp(43852) := x"6800";
    tmp(43853) := x"7000";
    tmp(43854) := x"7820";
    tmp(43855) := x"7820";
    tmp(43856) := x"8820";
    tmp(43857) := x"b821";
    tmp(43858) := x"d041";
    tmp(43859) := x"e861";
    tmp(43860) := x"6881";
    tmp(43861) := x"1040";
    tmp(43862) := x"0840";
    tmp(43863) := x"0840";
    tmp(43864) := x"0840";
    tmp(43865) := x"0840";
    tmp(43866) := x"0840";
    tmp(43867) := x"0840";
    tmp(43868) := x"0840";
    tmp(43869) := x"0840";
    tmp(43870) := x"0840";
    tmp(43871) := x"0840";
    tmp(43872) := x"0840";
    tmp(43873) := x"0840";
    tmp(43874) := x"0840";
    tmp(43875) := x"0840";
    tmp(43876) := x"0840";
    tmp(43877) := x"001f";
    tmp(43878) := x"001f";
    tmp(43879) := x"001f";
    tmp(43880) := x"001f";
    tmp(43881) := x"001f";
    tmp(43882) := x"001f";
    tmp(43883) := x"001f";
    tmp(43884) := x"001f";
    tmp(43885) := x"001f";
    tmp(43886) := x"001f";
    tmp(43887) := x"001f";
    tmp(43888) := x"001f";
    tmp(43889) := x"001f";
    tmp(43890) := x"001f";
    tmp(43891) := x"001f";
    tmp(43892) := x"001f";
    tmp(43893) := x"001f";
    tmp(43894) := x"001f";
    tmp(43895) := x"001f";
    tmp(43896) := x"001f";
    tmp(43897) := x"001f";
    tmp(43898) := x"001f";
    tmp(43899) := x"001f";
    tmp(43900) := x"001f";
    tmp(43901) := x"001f";
    tmp(43902) := x"001f";
    tmp(43903) := x"001f";
    tmp(43904) := x"001f";
    tmp(43905) := x"001f";
    tmp(43906) := x"001f";
    tmp(43907) := x"001f";
    tmp(43908) := x"001f";
    tmp(43909) := x"001f";
    tmp(43910) := x"001f";
    tmp(43911) := x"001f";
    tmp(43912) := x"001f";
    tmp(43913) := x"001f";
    tmp(43914) := x"001f";
    tmp(43915) := x"001f";
    tmp(43916) := x"001f";
    tmp(43917) := x"0840";
    tmp(43918) := x"1060";
    tmp(43919) := x"1061";
    tmp(43920) := x"0000";
    tmp(43921) := x"0880";
    tmp(43922) := x"0880";
    tmp(43923) := x"0880";
    tmp(43924) := x"0880";
    tmp(43925) := x"0880";
    tmp(43926) := x"0880";
    tmp(43927) := x"0880";
    tmp(43928) := x"0880";
    tmp(43929) := x"0880";
    tmp(43930) := x"0880";
    tmp(43931) := x"0880";
    tmp(43932) := x"0860";
    tmp(43933) := x"0860";
    tmp(43934) := x"0860";
    tmp(43935) := x"0860";
    tmp(43936) := x"0860";
    tmp(43937) := x"0840";
    tmp(43938) := x"0840";
    tmp(43939) := x"0840";
    tmp(43940) := x"0840";
    tmp(43941) := x"0840";
    tmp(43942) := x"0840";
    tmp(43943) := x"0840";
    tmp(43944) := x"0840";
    tmp(43945) := x"0840";
    tmp(43946) := x"0840";
    tmp(43947) := x"0840";
    tmp(43948) := x"0840";
    tmp(43949) := x"0840";
    tmp(43950) := x"0860";
    tmp(43951) := x"0860";
    tmp(43952) := x"0880";
    tmp(43953) := x"0880";
    tmp(43954) := x"0880";
    tmp(43955) := x"08a0";
    tmp(43956) := x"08a0";
    tmp(43957) := x"08a0";
    tmp(43958) := x"08a0";
    tmp(43959) := x"08a0";
    tmp(43960) := x"08a0";
    tmp(43961) := x"08c0";
    tmp(43962) := x"08c0";
    tmp(43963) := x"08e0";
    tmp(43964) := x"08e0";
    tmp(43965) := x"0900";
    tmp(43966) := x"0900";
    tmp(43967) := x"08e0";
    tmp(43968) := x"08e0";
    tmp(43969) := x"0900";
    tmp(43970) := x"0900";
    tmp(43971) := x"0900";
    tmp(43972) := x"0900";
    tmp(43973) := x"0900";
    tmp(43974) := x"0900";
    tmp(43975) := x"0900";
    tmp(43976) := x"0900";
    tmp(43977) := x"0920";
    tmp(43978) := x"0920";
    tmp(43979) := x"0920";
    tmp(43980) := x"0920";
    tmp(43981) := x"0920";
    tmp(43982) := x"0920";
    tmp(43983) := x"0920";
    tmp(43984) := x"0920";
    tmp(43985) := x"0900";
    tmp(43986) := x"0900";
    tmp(43987) := x"0900";
    tmp(43988) := x"0900";
    tmp(43989) := x"0900";
    tmp(43990) := x"0900";
    tmp(43991) := x"0900";
    tmp(43992) := x"0900";
    tmp(43993) := x"0900";
    tmp(43994) := x"0900";
    tmp(43995) := x"0900";
    tmp(43996) := x"08e0";
    tmp(43997) := x"08e0";
    tmp(43998) := x"08e0";
    tmp(43999) := x"08e0";
    tmp(44000) := x"08e0";
    tmp(44001) := x"08e0";
    tmp(44002) := x"08e0";
    tmp(44003) := x"08e0";
    tmp(44004) := x"08e0";
    tmp(44005) := x"0900";
    tmp(44006) := x"0900";
    tmp(44007) := x"0900";
    tmp(44008) := x"0900";
    tmp(44009) := x"0900";
    tmp(44010) := x"0900";
    tmp(44011) := x"0900";
    tmp(44012) := x"0900";
    tmp(44013) := x"0900";
    tmp(44014) := x"0920";
    tmp(44015) := x"0920";
    tmp(44016) := x"0920";
    tmp(44017) := x"0920";
    tmp(44018) := x"0920";
    tmp(44019) := x"0920";
    tmp(44020) := x"0920";
    tmp(44021) := x"0920";
    tmp(44022) := x"0900";
    tmp(44023) := x"0900";
    tmp(44024) := x"0900";
    tmp(44025) := x"08e0";
    tmp(44026) := x"08c0";
    tmp(44027) := x"2100";
    tmp(44028) := x"51a2";
    tmp(44029) := x"79e4";
    tmp(44030) := x"8225";
    tmp(44031) := x"8a46";
    tmp(44032) := x"9aa8";
    tmp(44033) := x"ab4c";
    tmp(44034) := x"b3ae";
    tmp(44035) := x"c410";
    tmp(44036) := x"c471";
    tmp(44037) := x"d472";
    tmp(44038) := x"cc30";
    tmp(44039) := x"cc30";
    tmp(44040) := x"c3cf";
    tmp(44041) := x"c38e";
    tmp(44042) := x"c36c";
    tmp(44043) := x"c38c";
    tmp(44044) := x"cbad";
    tmp(44045) := x"c34c";
    tmp(44046) := x"bb0b";
    tmp(44047) := x"b2ca";
    tmp(44048) := x"bb2b";
    tmp(44049) := x"c36c";
    tmp(44050) := x"bb2b";
    tmp(44051) := x"bb2a";
    tmp(44052) := x"d3cb";
    tmp(44053) := x"c34a";
    tmp(44054) := x"cb4a";
    tmp(44055) := x"bb08";
    tmp(44056) := x"c328";
    tmp(44057) := x"c349";
    tmp(44058) := x"cb8a";
    tmp(44059) := x"cb6a";
    tmp(44060) := x"b2e9";
    tmp(44061) := x"9a67";
    tmp(44062) := x"79c5";
    tmp(44063) := x"5944";
    tmp(44064) := x"4903";
    tmp(44065) := x"5985";
    tmp(44066) := x"4924";
    tmp(44067) := x"4944";
    tmp(44068) := x"4124";
    tmp(44069) := x"5165";
    tmp(44070) := x"5986";
    tmp(44071) := x"30e4";
    tmp(44072) := x"1862";
    tmp(44073) := x"1862";
    tmp(44074) := x"5104";
    tmp(44075) := x"89a6";
    tmp(44076) := x"7145";
    tmp(44077) := x"4082";
    tmp(44078) := x"1000";
    tmp(44079) := x"0800";
    tmp(44080) := x"1000";
    tmp(44081) := x"1000";
    tmp(44082) := x"1000";
    tmp(44083) := x"1000";
    tmp(44084) := x"1800";
    tmp(44085) := x"2000";
    tmp(44086) := x"3000";
    tmp(44087) := x"4000";
    tmp(44088) := x"4800";
    tmp(44089) := x"5000";
    tmp(44090) := x"5800";
    tmp(44091) := x"6000";
    tmp(44092) := x"6800";
    tmp(44093) := x"7800";
    tmp(44094) := x"8000";
    tmp(44095) := x"8820";
    tmp(44096) := x"8820";
    tmp(44097) := x"b020";
    tmp(44098) := x"b820";
    tmp(44099) := x"c821";
    tmp(44100) := x"b881";
    tmp(44101) := x"2840";
    tmp(44102) := x"1040";
    tmp(44103) := x"0840";
    tmp(44104) := x"0840";
    tmp(44105) := x"0840";
    tmp(44106) := x"0840";
    tmp(44107) := x"0840";
    tmp(44108) := x"0840";
    tmp(44109) := x"0840";
    tmp(44110) := x"0840";
    tmp(44111) := x"0840";
    tmp(44112) := x"0840";
    tmp(44113) := x"0840";
    tmp(44114) := x"0840";
    tmp(44115) := x"0840";
    tmp(44116) := x"0840";
    tmp(44117) := x"001f";
    tmp(44118) := x"001f";
    tmp(44119) := x"001f";
    tmp(44120) := x"001f";
    tmp(44121) := x"001f";
    tmp(44122) := x"001f";
    tmp(44123) := x"001f";
    tmp(44124) := x"001f";
    tmp(44125) := x"001f";
    tmp(44126) := x"001f";
    tmp(44127) := x"001f";
    tmp(44128) := x"001f";
    tmp(44129) := x"001f";
    tmp(44130) := x"001f";
    tmp(44131) := x"001f";
    tmp(44132) := x"001f";
    tmp(44133) := x"001f";
    tmp(44134) := x"001f";
    tmp(44135) := x"001f";
    tmp(44136) := x"001f";
    tmp(44137) := x"001f";
    tmp(44138) := x"001f";
    tmp(44139) := x"001f";
    tmp(44140) := x"001f";
    tmp(44141) := x"001f";
    tmp(44142) := x"001f";
    tmp(44143) := x"001f";
    tmp(44144) := x"001f";
    tmp(44145) := x"001f";
    tmp(44146) := x"001f";
    tmp(44147) := x"001f";
    tmp(44148) := x"001f";
    tmp(44149) := x"001f";
    tmp(44150) := x"001f";
    tmp(44151) := x"001f";
    tmp(44152) := x"001f";
    tmp(44153) := x"001f";
    tmp(44154) := x"001f";
    tmp(44155) := x"001f";
    tmp(44156) := x"001f";
    tmp(44157) := x"0840";
    tmp(44158) := x"1060";
    tmp(44159) := x"1060";
    tmp(44160) := x"0000";
    tmp(44161) := x"0880";
    tmp(44162) := x"0880";
    tmp(44163) := x"0880";
    tmp(44164) := x"0880";
    tmp(44165) := x"0880";
    tmp(44166) := x"0881";
    tmp(44167) := x"0880";
    tmp(44168) := x"0880";
    tmp(44169) := x"0880";
    tmp(44170) := x"0880";
    tmp(44171) := x"0880";
    tmp(44172) := x"0880";
    tmp(44173) := x"0880";
    tmp(44174) := x"0860";
    tmp(44175) := x"0860";
    tmp(44176) := x"0860";
    tmp(44177) := x"0860";
    tmp(44178) := x"0840";
    tmp(44179) := x"0840";
    tmp(44180) := x"0840";
    tmp(44181) := x"0840";
    tmp(44182) := x"0840";
    tmp(44183) := x"0840";
    tmp(44184) := x"0840";
    tmp(44185) := x"0840";
    tmp(44186) := x"0840";
    tmp(44187) := x"0840";
    tmp(44188) := x"0840";
    tmp(44189) := x"0840";
    tmp(44190) := x"0840";
    tmp(44191) := x"0860";
    tmp(44192) := x"0860";
    tmp(44193) := x"0860";
    tmp(44194) := x"0880";
    tmp(44195) := x"0880";
    tmp(44196) := x"0880";
    tmp(44197) := x"08a0";
    tmp(44198) := x"08a0";
    tmp(44199) := x"08a0";
    tmp(44200) := x"08a0";
    tmp(44201) := x"08a0";
    tmp(44202) := x"08c0";
    tmp(44203) := x"08c0";
    tmp(44204) := x"08c0";
    tmp(44205) := x"08e0";
    tmp(44206) := x"08e0";
    tmp(44207) := x"08e0";
    tmp(44208) := x"08e0";
    tmp(44209) := x"0900";
    tmp(44210) := x"0900";
    tmp(44211) := x"0900";
    tmp(44212) := x"0900";
    tmp(44213) := x"0900";
    tmp(44214) := x"0900";
    tmp(44215) := x"0900";
    tmp(44216) := x"0900";
    tmp(44217) := x"0900";
    tmp(44218) := x"0920";
    tmp(44219) := x"0900";
    tmp(44220) := x"0920";
    tmp(44221) := x"0920";
    tmp(44222) := x"0920";
    tmp(44223) := x"0920";
    tmp(44224) := x"0900";
    tmp(44225) := x"0900";
    tmp(44226) := x"0900";
    tmp(44227) := x"0900";
    tmp(44228) := x"0900";
    tmp(44229) := x"0900";
    tmp(44230) := x"0900";
    tmp(44231) := x"0900";
    tmp(44232) := x"0900";
    tmp(44233) := x"0900";
    tmp(44234) := x"0900";
    tmp(44235) := x"0900";
    tmp(44236) := x"08e0";
    tmp(44237) := x"08e0";
    tmp(44238) := x"08e0";
    tmp(44239) := x"08e0";
    tmp(44240) := x"08e0";
    tmp(44241) := x"08e0";
    tmp(44242) := x"08e0";
    tmp(44243) := x"08e0";
    tmp(44244) := x"08e0";
    tmp(44245) := x"0900";
    tmp(44246) := x"0900";
    tmp(44247) := x"0900";
    tmp(44248) := x"0900";
    tmp(44249) := x"0900";
    tmp(44250) := x"0920";
    tmp(44251) := x"0920";
    tmp(44252) := x"0900";
    tmp(44253) := x"0920";
    tmp(44254) := x"0920";
    tmp(44255) := x"0920";
    tmp(44256) := x"0920";
    tmp(44257) := x"0920";
    tmp(44258) := x"0920";
    tmp(44259) := x"0920";
    tmp(44260) := x"0920";
    tmp(44261) := x"0920";
    tmp(44262) := x"0900";
    tmp(44263) := x"0900";
    tmp(44264) := x"0900";
    tmp(44265) := x"08c0";
    tmp(44266) := x"2141";
    tmp(44267) := x"51a2";
    tmp(44268) := x"71e4";
    tmp(44269) := x"8225";
    tmp(44270) := x"8a67";
    tmp(44271) := x"9aea";
    tmp(44272) := x"ab4c";
    tmp(44273) := x"ab6d";
    tmp(44274) := x"b38e";
    tmp(44275) := x"bbef";
    tmp(44276) := x"bc0f";
    tmp(44277) := x"c3ef";
    tmp(44278) := x"c3ce";
    tmp(44279) := x"c3ce";
    tmp(44280) := x"bb8e";
    tmp(44281) := x"bb6d";
    tmp(44282) := x"bb2b";
    tmp(44283) := x"bb4c";
    tmp(44284) := x"c38d";
    tmp(44285) := x"c38d";
    tmp(44286) := x"b32b";
    tmp(44287) := x"aac9";
    tmp(44288) := x"b30a";
    tmp(44289) := x"bb2b";
    tmp(44290) := x"bb0a";
    tmp(44291) := x"bb2a";
    tmp(44292) := x"bb4a";
    tmp(44293) := x"c34a";
    tmp(44294) := x"c349";
    tmp(44295) := x"bb08";
    tmp(44296) := x"c328";
    tmp(44297) := x"bb09";
    tmp(44298) := x"cbab";
    tmp(44299) := x"cbac";
    tmp(44300) := x"aae9";
    tmp(44301) := x"b309";
    tmp(44302) := x"9267";
    tmp(44303) := x"5144";
    tmp(44304) := x"30a2";
    tmp(44305) := x"30a2";
    tmp(44306) := x"1861";
    tmp(44307) := x"1861";
    tmp(44308) := x"1061";
    tmp(44309) := x"2082";
    tmp(44310) := x"20a2";
    tmp(44311) := x"20a3";
    tmp(44312) := x"20c4";
    tmp(44313) := x"20a2";
    tmp(44314) := x"71a6";
    tmp(44315) := x"6925";
    tmp(44316) := x"6104";
    tmp(44317) := x"2041";
    tmp(44318) := x"0800";
    tmp(44319) := x"0800";
    tmp(44320) := x"1000";
    tmp(44321) := x"1000";
    tmp(44322) := x"1000";
    tmp(44323) := x"1800";
    tmp(44324) := x"1800";
    tmp(44325) := x"2800";
    tmp(44326) := x"3000";
    tmp(44327) := x"3800";
    tmp(44328) := x"4000";
    tmp(44329) := x"5000";
    tmp(44330) := x"5800";
    tmp(44331) := x"6000";
    tmp(44332) := x"6800";
    tmp(44333) := x"7000";
    tmp(44334) := x"8800";
    tmp(44335) := x"9820";
    tmp(44336) := x"a020";
    tmp(44337) := x"a820";
    tmp(44338) := x"c821";
    tmp(44339) := x"d041";
    tmp(44340) := x"e041";
    tmp(44341) := x"7861";
    tmp(44342) := x"1040";
    tmp(44343) := x"1040";
    tmp(44344) := x"0840";
    tmp(44345) := x"0840";
    tmp(44346) := x"0840";
    tmp(44347) := x"0840";
    tmp(44348) := x"0840";
    tmp(44349) := x"0840";
    tmp(44350) := x"0840";
    tmp(44351) := x"0840";
    tmp(44352) := x"0840";
    tmp(44353) := x"0840";
    tmp(44354) := x"0840";
    tmp(44355) := x"0840";
    tmp(44356) := x"0840";
    tmp(44357) := x"001f";
    tmp(44358) := x"001f";
    tmp(44359) := x"001f";
    tmp(44360) := x"001f";
    tmp(44361) := x"001f";
    tmp(44362) := x"001f";
    tmp(44363) := x"001f";
    tmp(44364) := x"001f";
    tmp(44365) := x"001f";
    tmp(44366) := x"001f";
    tmp(44367) := x"001f";
    tmp(44368) := x"001f";
    tmp(44369) := x"001f";
    tmp(44370) := x"001f";
    tmp(44371) := x"001f";
    tmp(44372) := x"001f";
    tmp(44373) := x"001f";
    tmp(44374) := x"001f";
    tmp(44375) := x"001f";
    tmp(44376) := x"001f";
    tmp(44377) := x"001f";
    tmp(44378) := x"001f";
    tmp(44379) := x"001f";
    tmp(44380) := x"001f";
    tmp(44381) := x"001f";
    tmp(44382) := x"001f";
    tmp(44383) := x"001f";
    tmp(44384) := x"001f";
    tmp(44385) := x"001f";
    tmp(44386) := x"001f";
    tmp(44387) := x"001f";
    tmp(44388) := x"001f";
    tmp(44389) := x"001f";
    tmp(44390) := x"001f";
    tmp(44391) := x"001f";
    tmp(44392) := x"001f";
    tmp(44393) := x"001f";
    tmp(44394) := x"001f";
    tmp(44395) := x"001f";
    tmp(44396) := x"001f";
    tmp(44397) := x"0840";
    tmp(44398) := x"1061";
    tmp(44399) := x"0860";
    tmp(44400) := x"0000";
    tmp(44401) := x"08a0";
    tmp(44402) := x"08a0";
    tmp(44403) := x"0881";
    tmp(44404) := x"0881";
    tmp(44405) := x"0881";
    tmp(44406) := x"0881";
    tmp(44407) := x"0881";
    tmp(44408) := x"0881";
    tmp(44409) := x"0881";
    tmp(44410) := x"0881";
    tmp(44411) := x"0880";
    tmp(44412) := x"0880";
    tmp(44413) := x"0880";
    tmp(44414) := x"0880";
    tmp(44415) := x"0860";
    tmp(44416) := x"0860";
    tmp(44417) := x"0860";
    tmp(44418) := x"0860";
    tmp(44419) := x"0840";
    tmp(44420) := x"0840";
    tmp(44421) := x"0840";
    tmp(44422) := x"0840";
    tmp(44423) := x"0840";
    tmp(44424) := x"0840";
    tmp(44425) := x"0840";
    tmp(44426) := x"0840";
    tmp(44427) := x"0840";
    tmp(44428) := x"0840";
    tmp(44429) := x"0840";
    tmp(44430) := x"0840";
    tmp(44431) := x"0860";
    tmp(44432) := x"0860";
    tmp(44433) := x"0860";
    tmp(44434) := x"0860";
    tmp(44435) := x"0880";
    tmp(44436) := x"0880";
    tmp(44437) := x"0880";
    tmp(44438) := x"0880";
    tmp(44439) := x"0880";
    tmp(44440) := x"08a0";
    tmp(44441) := x"08a0";
    tmp(44442) := x"08a0";
    tmp(44443) := x"08c0";
    tmp(44444) := x"08c0";
    tmp(44445) := x"08c0";
    tmp(44446) := x"08c0";
    tmp(44447) := x"08e0";
    tmp(44448) := x"08e0";
    tmp(44449) := x"08e0";
    tmp(44450) := x"0900";
    tmp(44451) := x"08e0";
    tmp(44452) := x"0900";
    tmp(44453) := x"0900";
    tmp(44454) := x"0900";
    tmp(44455) := x"0900";
    tmp(44456) := x"0900";
    tmp(44457) := x"0920";
    tmp(44458) := x"0900";
    tmp(44459) := x"0900";
    tmp(44460) := x"0920";
    tmp(44461) := x"0900";
    tmp(44462) := x"0900";
    tmp(44463) := x"0920";
    tmp(44464) := x"0900";
    tmp(44465) := x"0900";
    tmp(44466) := x"0900";
    tmp(44467) := x"0900";
    tmp(44468) := x"0900";
    tmp(44469) := x"0900";
    tmp(44470) := x"0900";
    tmp(44471) := x"0900";
    tmp(44472) := x"0900";
    tmp(44473) := x"0900";
    tmp(44474) := x"0900";
    tmp(44475) := x"08e0";
    tmp(44476) := x"08e0";
    tmp(44477) := x"08e0";
    tmp(44478) := x"08e0";
    tmp(44479) := x"08e0";
    tmp(44480) := x"08e0";
    tmp(44481) := x"08e0";
    tmp(44482) := x"0900";
    tmp(44483) := x"0900";
    tmp(44484) := x"08e0";
    tmp(44485) := x"0900";
    tmp(44486) := x"0900";
    tmp(44487) := x"0900";
    tmp(44488) := x"0900";
    tmp(44489) := x"0900";
    tmp(44490) := x"0900";
    tmp(44491) := x"0900";
    tmp(44492) := x"0920";
    tmp(44493) := x"0920";
    tmp(44494) := x"0920";
    tmp(44495) := x"0920";
    tmp(44496) := x"0920";
    tmp(44497) := x"0920";
    tmp(44498) := x"0920";
    tmp(44499) := x"0920";
    tmp(44500) := x"0920";
    tmp(44501) := x"0920";
    tmp(44502) := x"0920";
    tmp(44503) := x"0900";
    tmp(44504) := x"08c0";
    tmp(44505) := x"1920";
    tmp(44506) := x"51a2";
    tmp(44507) := x"69e4";
    tmp(44508) := x"7a25";
    tmp(44509) := x"92a8";
    tmp(44510) := x"a32b";
    tmp(44511) := x"a36d";
    tmp(44512) := x"a36d";
    tmp(44513) := x"ab8d";
    tmp(44514) := x"b36d";
    tmp(44515) := x"bbce";
    tmp(44516) := x"bbce";
    tmp(44517) := x"bbae";
    tmp(44518) := x"bb8d";
    tmp(44519) := x"ab4b";
    tmp(44520) := x"ab2b";
    tmp(44521) := x"b32b";
    tmp(44522) := x"b2eb";
    tmp(44523) := x"b30b";
    tmp(44524) := x"b32c";
    tmp(44525) := x"bb8d";
    tmp(44526) := x"b34c";
    tmp(44527) := x"b2ea";
    tmp(44528) := x"bb4b";
    tmp(44529) := x"b32b";
    tmp(44530) := x"b30a";
    tmp(44531) := x"bb2a";
    tmp(44532) := x"bb29";
    tmp(44533) := x"bb09";
    tmp(44534) := x"b308";
    tmp(44535) := x"c349";
    tmp(44536) := x"c349";
    tmp(44537) := x"bb29";
    tmp(44538) := x"cbab";
    tmp(44539) := x"cbed";
    tmp(44540) := x"c38c";
    tmp(44541) := x"dc0d";
    tmp(44542) := x"bb6b";
    tmp(44543) := x"9ac9";
    tmp(44544) := x"7206";
    tmp(44545) := x"5165";
    tmp(44546) := x"28a2";
    tmp(44547) := x"1861";
    tmp(44548) := x"1041";
    tmp(44549) := x"1041";
    tmp(44550) := x"1062";
    tmp(44551) := x"18c3";
    tmp(44552) := x"3125";
    tmp(44553) := x"30e3";
    tmp(44554) := x"8a07";
    tmp(44555) := x"60e4";
    tmp(44556) := x"48a2";
    tmp(44557) := x"0800";
    tmp(44558) := x"0800";
    tmp(44559) := x"1000";
    tmp(44560) := x"1000";
    tmp(44561) := x"1000";
    tmp(44562) := x"1000";
    tmp(44563) := x"2000";
    tmp(44564) := x"2000";
    tmp(44565) := x"2800";
    tmp(44566) := x"3000";
    tmp(44567) := x"3800";
    tmp(44568) := x"4000";
    tmp(44569) := x"5000";
    tmp(44570) := x"5800";
    tmp(44571) := x"6800";
    tmp(44572) := x"6800";
    tmp(44573) := x"6800";
    tmp(44574) := x"7800";
    tmp(44575) := x"9000";
    tmp(44576) := x"a020";
    tmp(44577) := x"b020";
    tmp(44578) := x"b820";
    tmp(44579) := x"d021";
    tmp(44580) := x"b820";
    tmp(44581) := x"c041";
    tmp(44582) := x"3861";
    tmp(44583) := x"1040";
    tmp(44584) := x"1040";
    tmp(44585) := x"0840";
    tmp(44586) := x"0840";
    tmp(44587) := x"0840";
    tmp(44588) := x"0840";
    tmp(44589) := x"0840";
    tmp(44590) := x"0840";
    tmp(44591) := x"0840";
    tmp(44592) := x"0840";
    tmp(44593) := x"0840";
    tmp(44594) := x"0840";
    tmp(44595) := x"0840";
    tmp(44596) := x"0840";
    tmp(44597) := x"001f";
    tmp(44598) := x"001f";
    tmp(44599) := x"001f";
    tmp(44600) := x"001f";
    tmp(44601) := x"001f";
    tmp(44602) := x"001f";
    tmp(44603) := x"001f";
    tmp(44604) := x"001f";
    tmp(44605) := x"001f";
    tmp(44606) := x"001f";
    tmp(44607) := x"001f";
    tmp(44608) := x"001f";
    tmp(44609) := x"001f";
    tmp(44610) := x"001f";
    tmp(44611) := x"001f";
    tmp(44612) := x"001f";
    tmp(44613) := x"001f";
    tmp(44614) := x"001f";
    tmp(44615) := x"001f";
    tmp(44616) := x"001f";
    tmp(44617) := x"001f";
    tmp(44618) := x"001f";
    tmp(44619) := x"001f";
    tmp(44620) := x"001f";
    tmp(44621) := x"001f";
    tmp(44622) := x"001f";
    tmp(44623) := x"001f";
    tmp(44624) := x"001f";
    tmp(44625) := x"001f";
    tmp(44626) := x"001f";
    tmp(44627) := x"001f";
    tmp(44628) := x"001f";
    tmp(44629) := x"001f";
    tmp(44630) := x"001f";
    tmp(44631) := x"001f";
    tmp(44632) := x"001f";
    tmp(44633) := x"001f";
    tmp(44634) := x"001f";
    tmp(44635) := x"001f";
    tmp(44636) := x"001f";
    tmp(44637) := x"0840";
    tmp(44638) := x"0840";
    tmp(44639) := x"0840";
    tmp(44640) := x"0000";
    tmp(44641) := x"08a0";
    tmp(44642) := x"0880";
    tmp(44643) := x"08a1";
    tmp(44644) := x"08a1";
    tmp(44645) := x"08a1";
    tmp(44646) := x"0881";
    tmp(44647) := x"08a1";
    tmp(44648) := x"08a1";
    tmp(44649) := x"0881";
    tmp(44650) := x"0881";
    tmp(44651) := x"0881";
    tmp(44652) := x"0881";
    tmp(44653) := x"0881";
    tmp(44654) := x"0881";
    tmp(44655) := x"0881";
    tmp(44656) := x"0880";
    tmp(44657) := x"0860";
    tmp(44658) := x"0860";
    tmp(44659) := x"0860";
    tmp(44660) := x"0840";
    tmp(44661) := x"0840";
    tmp(44662) := x"0840";
    tmp(44663) := x"0840";
    tmp(44664) := x"0840";
    tmp(44665) := x"0840";
    tmp(44666) := x"0840";
    tmp(44667) := x"0840";
    tmp(44668) := x"0840";
    tmp(44669) := x"0840";
    tmp(44670) := x"0840";
    tmp(44671) := x"0840";
    tmp(44672) := x"0860";
    tmp(44673) := x"0860";
    tmp(44674) := x"0860";
    tmp(44675) := x"0860";
    tmp(44676) := x"0860";
    tmp(44677) := x"0880";
    tmp(44678) := x"0880";
    tmp(44679) := x"0880";
    tmp(44680) := x"0880";
    tmp(44681) := x"0880";
    tmp(44682) := x"08a0";
    tmp(44683) := x"08a0";
    tmp(44684) := x"08a0";
    tmp(44685) := x"08c0";
    tmp(44686) := x"08c0";
    tmp(44687) := x"08e0";
    tmp(44688) := x"08e0";
    tmp(44689) := x"08e0";
    tmp(44690) := x"08e0";
    tmp(44691) := x"08e0";
    tmp(44692) := x"0900";
    tmp(44693) := x"0900";
    tmp(44694) := x"0900";
    tmp(44695) := x"0900";
    tmp(44696) := x"0900";
    tmp(44697) := x"0900";
    tmp(44698) := x"0900";
    tmp(44699) := x"0900";
    tmp(44700) := x"0920";
    tmp(44701) := x"0900";
    tmp(44702) := x"0920";
    tmp(44703) := x"0900";
    tmp(44704) := x"0920";
    tmp(44705) := x"0920";
    tmp(44706) := x"0900";
    tmp(44707) := x"0900";
    tmp(44708) := x"0900";
    tmp(44709) := x"0900";
    tmp(44710) := x"0900";
    tmp(44711) := x"0900";
    tmp(44712) := x"0900";
    tmp(44713) := x"0900";
    tmp(44714) := x"0900";
    tmp(44715) := x"0900";
    tmp(44716) := x"08e0";
    tmp(44717) := x"08e0";
    tmp(44718) := x"08e0";
    tmp(44719) := x"08e0";
    tmp(44720) := x"08e0";
    tmp(44721) := x"08e0";
    tmp(44722) := x"08e0";
    tmp(44723) := x"0900";
    tmp(44724) := x"0900";
    tmp(44725) := x"0900";
    tmp(44726) := x"0900";
    tmp(44727) := x"0900";
    tmp(44728) := x"0900";
    tmp(44729) := x"0900";
    tmp(44730) := x"0900";
    tmp(44731) := x"0920";
    tmp(44732) := x"0920";
    tmp(44733) := x"0920";
    tmp(44734) := x"0920";
    tmp(44735) := x"0920";
    tmp(44736) := x"0920";
    tmp(44737) := x"0920";
    tmp(44738) := x"0920";
    tmp(44739) := x"0920";
    tmp(44740) := x"0920";
    tmp(44741) := x"0920";
    tmp(44742) := x"0900";
    tmp(44743) := x"0900";
    tmp(44744) := x"10e0";
    tmp(44745) := x"49a2";
    tmp(44746) := x"6a04";
    tmp(44747) := x"7a46";
    tmp(44748) := x"92e9";
    tmp(44749) := x"ab6d";
    tmp(44750) := x"abae";
    tmp(44751) := x"ab8e";
    tmp(44752) := x"a36d";
    tmp(44753) := x"ab8e";
    tmp(44754) := x"ab8e";
    tmp(44755) := x"bbef";
    tmp(44756) := x"bbcf";
    tmp(44757) := x"b3ae";
    tmp(44758) := x"ab4c";
    tmp(44759) := x"9aca";
    tmp(44760) := x"9289";
    tmp(44761) := x"ab2b";
    tmp(44762) := x"b30b";
    tmp(44763) := x"aaeb";
    tmp(44764) := x"ab0b";
    tmp(44765) := x"b34c";
    tmp(44766) := x"b34d";
    tmp(44767) := x"a2ca";
    tmp(44768) := x"aaea";
    tmp(44769) := x"bb4c";
    tmp(44770) := x"bb4b";
    tmp(44771) := x"b30a";
    tmp(44772) := x"b309";
    tmp(44773) := x"b2e9";
    tmp(44774) := x"b309";
    tmp(44775) := x"c38a";
    tmp(44776) := x"bb29";
    tmp(44777) := x"c34a";
    tmp(44778) := x"bb4a";
    tmp(44779) := x"c3cc";
    tmp(44780) := x"cbcd";
    tmp(44781) := x"bb6b";
    tmp(44782) := x"cbac";
    tmp(44783) := x"c3ed";
    tmp(44784) := x"b34b";
    tmp(44785) := x"ab4b";
    tmp(44786) := x"8a89";
    tmp(44787) := x"5186";
    tmp(44788) := x"20a2";
    tmp(44789) := x"1882";
    tmp(44790) := x"1041";
    tmp(44791) := x"1062";
    tmp(44792) := x"20a3";
    tmp(44793) := x"5985";
    tmp(44794) := x"7144";
    tmp(44795) := x"4061";
    tmp(44796) := x"2020";
    tmp(44797) := x"0800";
    tmp(44798) := x"1000";
    tmp(44799) := x"1000";
    tmp(44800) := x"1000";
    tmp(44801) := x"1000";
    tmp(44802) := x"1000";
    tmp(44803) := x"1800";
    tmp(44804) := x"2000";
    tmp(44805) := x"2800";
    tmp(44806) := x"3800";
    tmp(44807) := x"4000";
    tmp(44808) := x"4800";
    tmp(44809) := x"5800";
    tmp(44810) := x"6000";
    tmp(44811) := x"7000";
    tmp(44812) := x"7820";
    tmp(44813) := x"6800";
    tmp(44814) := x"7000";
    tmp(44815) := x"8800";
    tmp(44816) := x"a020";
    tmp(44817) := x"9800";
    tmp(44818) := x"c020";
    tmp(44819) := x"c020";
    tmp(44820) := x"a820";
    tmp(44821) := x"b820";
    tmp(44822) := x"6061";
    tmp(44823) := x"1040";
    tmp(44824) := x"1040";
    tmp(44825) := x"0840";
    tmp(44826) := x"0840";
    tmp(44827) := x"0840";
    tmp(44828) := x"0840";
    tmp(44829) := x"0840";
    tmp(44830) := x"0840";
    tmp(44831) := x"0840";
    tmp(44832) := x"0840";
    tmp(44833) := x"0840";
    tmp(44834) := x"0840";
    tmp(44835) := x"0840";
    tmp(44836) := x"0840";
    tmp(44837) := x"001f";
    tmp(44838) := x"001f";
    tmp(44839) := x"001f";
    tmp(44840) := x"001f";
    tmp(44841) := x"001f";
    tmp(44842) := x"001f";
    tmp(44843) := x"001f";
    tmp(44844) := x"001f";
    tmp(44845) := x"001f";
    tmp(44846) := x"001f";
    tmp(44847) := x"001f";
    tmp(44848) := x"001f";
    tmp(44849) := x"001f";
    tmp(44850) := x"001f";
    tmp(44851) := x"001f";
    tmp(44852) := x"001f";
    tmp(44853) := x"001f";
    tmp(44854) := x"001f";
    tmp(44855) := x"001f";
    tmp(44856) := x"001f";
    tmp(44857) := x"001f";
    tmp(44858) := x"001f";
    tmp(44859) := x"001f";
    tmp(44860) := x"001f";
    tmp(44861) := x"001f";
    tmp(44862) := x"001f";
    tmp(44863) := x"001f";
    tmp(44864) := x"001f";
    tmp(44865) := x"001f";
    tmp(44866) := x"001f";
    tmp(44867) := x"001f";
    tmp(44868) := x"001f";
    tmp(44869) := x"001f";
    tmp(44870) := x"001f";
    tmp(44871) := x"001f";
    tmp(44872) := x"001f";
    tmp(44873) := x"001f";
    tmp(44874) := x"001f";
    tmp(44875) := x"001f";
    tmp(44876) := x"001f";
    tmp(44877) := x"0840";
    tmp(44878) := x"0840";
    tmp(44879) := x"0840";
    tmp(44880) := x"0000";
    tmp(44881) := x"08a1";
    tmp(44882) := x"0880";
    tmp(44883) := x"08a0";
    tmp(44884) := x"08a1";
    tmp(44885) := x"08a1";
    tmp(44886) := x"08a1";
    tmp(44887) := x"08a1";
    tmp(44888) := x"08a1";
    tmp(44889) := x"0881";
    tmp(44890) := x"08a1";
    tmp(44891) := x"08a1";
    tmp(44892) := x"1081";
    tmp(44893) := x"0881";
    tmp(44894) := x"0881";
    tmp(44895) := x"0881";
    tmp(44896) := x"0881";
    tmp(44897) := x"0880";
    tmp(44898) := x"0860";
    tmp(44899) := x"0860";
    tmp(44900) := x"0860";
    tmp(44901) := x"0860";
    tmp(44902) := x"0840";
    tmp(44903) := x"0840";
    tmp(44904) := x"0840";
    tmp(44905) := x"0840";
    tmp(44906) := x"0840";
    tmp(44907) := x"0840";
    tmp(44908) := x"0840";
    tmp(44909) := x"0840";
    tmp(44910) := x"0840";
    tmp(44911) := x"0840";
    tmp(44912) := x"0860";
    tmp(44913) := x"0860";
    tmp(44914) := x"0860";
    tmp(44915) := x"0860";
    tmp(44916) := x"0860";
    tmp(44917) := x"0860";
    tmp(44918) := x"0860";
    tmp(44919) := x"0880";
    tmp(44920) := x"0880";
    tmp(44921) := x"0880";
    tmp(44922) := x"0880";
    tmp(44923) := x"0880";
    tmp(44924) := x"08a0";
    tmp(44925) := x"08a0";
    tmp(44926) := x"08c0";
    tmp(44927) := x"08c0";
    tmp(44928) := x"08c0";
    tmp(44929) := x"08e0";
    tmp(44930) := x"08e0";
    tmp(44931) := x"08e0";
    tmp(44932) := x"08e0";
    tmp(44933) := x"08e0";
    tmp(44934) := x"0900";
    tmp(44935) := x"0900";
    tmp(44936) := x"08e0";
    tmp(44937) := x"0900";
    tmp(44938) := x"0920";
    tmp(44939) := x"0920";
    tmp(44940) := x"0920";
    tmp(44941) := x"0920";
    tmp(44942) := x"0920";
    tmp(44943) := x"0920";
    tmp(44944) := x"0920";
    tmp(44945) := x"0900";
    tmp(44946) := x"0920";
    tmp(44947) := x"0900";
    tmp(44948) := x"0900";
    tmp(44949) := x"0900";
    tmp(44950) := x"0900";
    tmp(44951) := x"0900";
    tmp(44952) := x"0900";
    tmp(44953) := x"0900";
    tmp(44954) := x"08e0";
    tmp(44955) := x"0900";
    tmp(44956) := x"08e0";
    tmp(44957) := x"08e0";
    tmp(44958) := x"08e0";
    tmp(44959) := x"08e0";
    tmp(44960) := x"08e0";
    tmp(44961) := x"08e0";
    tmp(44962) := x"08e0";
    tmp(44963) := x"0900";
    tmp(44964) := x"0900";
    tmp(44965) := x"0900";
    tmp(44966) := x"0900";
    tmp(44967) := x"0900";
    tmp(44968) := x"0900";
    tmp(44969) := x"0900";
    tmp(44970) := x"0920";
    tmp(44971) := x"0920";
    tmp(44972) := x"0920";
    tmp(44973) := x"0920";
    tmp(44974) := x"0920";
    tmp(44975) := x"0920";
    tmp(44976) := x"0940";
    tmp(44977) := x"0920";
    tmp(44978) := x"0920";
    tmp(44979) := x"0920";
    tmp(44980) := x"0920";
    tmp(44981) := x"0920";
    tmp(44982) := x"0900";
    tmp(44983) := x"10e0";
    tmp(44984) := x"3161";
    tmp(44985) := x"61e4";
    tmp(44986) := x"7a67";
    tmp(44987) := x"92ea";
    tmp(44988) := x"9b4c";
    tmp(44989) := x"abae";
    tmp(44990) := x"a3af";
    tmp(44991) := x"9b8e";
    tmp(44992) := x"a3ae";
    tmp(44993) := x"b410";
    tmp(44994) := x"b3cf";
    tmp(44995) := x"a38e";
    tmp(44996) := x"abce";
    tmp(44997) := x"abae";
    tmp(44998) := x"a34d";
    tmp(44999) := x"9aeb";
    tmp(45000) := x"a2eb";
    tmp(45001) := x"9aca";
    tmp(45002) := x"a2ea";
    tmp(45003) := x"a30b";
    tmp(45004) := x"ab6d";
    tmp(45005) := x"a30b";
    tmp(45006) := x"92ca";
    tmp(45007) := x"8a68";
    tmp(45008) := x"9aa9";
    tmp(45009) := x"a30b";
    tmp(45010) := x"a2ca";
    tmp(45011) := x"b30a";
    tmp(45012) := x"aac8";
    tmp(45013) := x"b2e9";
    tmp(45014) := x"aae9";
    tmp(45015) := x"b329";
    tmp(45016) := x"b309";
    tmp(45017) := x"b30a";
    tmp(45018) := x"b30a";
    tmp(45019) := x"c3ac";
    tmp(45020) := x"bb4b";
    tmp(45021) := x"bb6b";
    tmp(45022) := x"c36b";
    tmp(45023) := x"c3ad";
    tmp(45024) := x"c3ce";
    tmp(45025) := x"b36d";
    tmp(45026) := x"a34c";
    tmp(45027) := x"7227";
    tmp(45028) := x"30e3";
    tmp(45029) := x"20a2";
    tmp(45030) := x"2904";
    tmp(45031) := x"20a2";
    tmp(45032) := x"2082";
    tmp(45033) := x"5103";
    tmp(45034) := x"3841";
    tmp(45035) := x"1800";
    tmp(45036) := x"1800";
    tmp(45037) := x"2000";
    tmp(45038) := x"3041";
    tmp(45039) := x"2020";
    tmp(45040) := x"1000";
    tmp(45041) := x"1800";
    tmp(45042) := x"1000";
    tmp(45043) := x"1000";
    tmp(45044) := x"1800";
    tmp(45045) := x"2800";
    tmp(45046) := x"3800";
    tmp(45047) := x"4800";
    tmp(45048) := x"5000";
    tmp(45049) := x"5800";
    tmp(45050) := x"6000";
    tmp(45051) := x"6800";
    tmp(45052) := x"7000";
    tmp(45053) := x"7800";
    tmp(45054) := x"7800";
    tmp(45055) := x"9000";
    tmp(45056) := x"a020";
    tmp(45057) := x"a820";
    tmp(45058) := x"c020";
    tmp(45059) := x"b020";
    tmp(45060) := x"c020";
    tmp(45061) := x"c020";
    tmp(45062) := x"9061";
    tmp(45063) := x"1840";
    tmp(45064) := x"1040";
    tmp(45065) := x"1040";
    tmp(45066) := x"0840";
    tmp(45067) := x"0840";
    tmp(45068) := x"0840";
    tmp(45069) := x"0840";
    tmp(45070) := x"0840";
    tmp(45071) := x"0840";
    tmp(45072) := x"0840";
    tmp(45073) := x"0840";
    tmp(45074) := x"0840";
    tmp(45075) := x"0840";
    tmp(45076) := x"0840";
    tmp(45077) := x"001f";
    tmp(45078) := x"001f";
    tmp(45079) := x"001f";
    tmp(45080) := x"001f";
    tmp(45081) := x"001f";
    tmp(45082) := x"001f";
    tmp(45083) := x"001f";
    tmp(45084) := x"001f";
    tmp(45085) := x"001f";
    tmp(45086) := x"001f";
    tmp(45087) := x"001f";
    tmp(45088) := x"001f";
    tmp(45089) := x"001f";
    tmp(45090) := x"001f";
    tmp(45091) := x"001f";
    tmp(45092) := x"001f";
    tmp(45093) := x"001f";
    tmp(45094) := x"001f";
    tmp(45095) := x"001f";
    tmp(45096) := x"001f";
    tmp(45097) := x"001f";
    tmp(45098) := x"001f";
    tmp(45099) := x"001f";
    tmp(45100) := x"001f";
    tmp(45101) := x"001f";
    tmp(45102) := x"001f";
    tmp(45103) := x"001f";
    tmp(45104) := x"001f";
    tmp(45105) := x"001f";
    tmp(45106) := x"001f";
    tmp(45107) := x"001f";
    tmp(45108) := x"001f";
    tmp(45109) := x"001f";
    tmp(45110) := x"001f";
    tmp(45111) := x"001f";
    tmp(45112) := x"001f";
    tmp(45113) := x"001f";
    tmp(45114) := x"001f";
    tmp(45115) := x"001f";
    tmp(45116) := x"001f";
    tmp(45117) := x"0840";
    tmp(45118) := x"0840";
    tmp(45119) := x"0840";
    tmp(45120) := x"0000";
    tmp(45121) := x"08a1";
    tmp(45122) := x"08a1";
    tmp(45123) := x"08a1";
    tmp(45124) := x"08a1";
    tmp(45125) := x"08a1";
    tmp(45126) := x"08a1";
    tmp(45127) := x"08a1";
    tmp(45128) := x"08a1";
    tmp(45129) := x"08a1";
    tmp(45130) := x"08a1";
    tmp(45131) := x"08a1";
    tmp(45132) := x"0881";
    tmp(45133) := x"10a1";
    tmp(45134) := x"10a1";
    tmp(45135) := x"0881";
    tmp(45136) := x"0881";
    tmp(45137) := x"0881";
    tmp(45138) := x"0881";
    tmp(45139) := x"0860";
    tmp(45140) := x"0860";
    tmp(45141) := x"0860";
    tmp(45142) := x"0860";
    tmp(45143) := x"0860";
    tmp(45144) := x"0860";
    tmp(45145) := x"0840";
    tmp(45146) := x"0840";
    tmp(45147) := x"0860";
    tmp(45148) := x"0860";
    tmp(45149) := x"0860";
    tmp(45150) := x"0860";
    tmp(45151) := x"0860";
    tmp(45152) := x"0840";
    tmp(45153) := x"0860";
    tmp(45154) := x"0860";
    tmp(45155) := x"0860";
    tmp(45156) := x"0860";
    tmp(45157) := x"0860";
    tmp(45158) := x"0860";
    tmp(45159) := x"0860";
    tmp(45160) := x"0860";
    tmp(45161) := x"0880";
    tmp(45162) := x"0880";
    tmp(45163) := x"0880";
    tmp(45164) := x"0880";
    tmp(45165) := x"08a0";
    tmp(45166) := x"08a0";
    tmp(45167) := x"08a0";
    tmp(45168) := x"08c0";
    tmp(45169) := x"08c0";
    tmp(45170) := x"08c0";
    tmp(45171) := x"08e0";
    tmp(45172) := x"08e0";
    tmp(45173) := x"08e0";
    tmp(45174) := x"08e0";
    tmp(45175) := x"08e0";
    tmp(45176) := x"0900";
    tmp(45177) := x"0900";
    tmp(45178) := x"0900";
    tmp(45179) := x"0920";
    tmp(45180) := x"0920";
    tmp(45181) := x"0920";
    tmp(45182) := x"0920";
    tmp(45183) := x"0920";
    tmp(45184) := x"0900";
    tmp(45185) := x"0900";
    tmp(45186) := x"0920";
    tmp(45187) := x"0900";
    tmp(45188) := x"0900";
    tmp(45189) := x"0920";
    tmp(45190) := x"0900";
    tmp(45191) := x"0900";
    tmp(45192) := x"0900";
    tmp(45193) := x"0900";
    tmp(45194) := x"08e0";
    tmp(45195) := x"08e0";
    tmp(45196) := x"0900";
    tmp(45197) := x"08e0";
    tmp(45198) := x"08e0";
    tmp(45199) := x"08e0";
    tmp(45200) := x"08e0";
    tmp(45201) := x"0900";
    tmp(45202) := x"0900";
    tmp(45203) := x"0900";
    tmp(45204) := x"0900";
    tmp(45205) := x"0900";
    tmp(45206) := x"0900";
    tmp(45207) := x"0900";
    tmp(45208) := x"0900";
    tmp(45209) := x"0920";
    tmp(45210) := x"0920";
    tmp(45211) := x"0920";
    tmp(45212) := x"0920";
    tmp(45213) := x"0920";
    tmp(45214) := x"0920";
    tmp(45215) := x"0920";
    tmp(45216) := x"0920";
    tmp(45217) := x"0920";
    tmp(45218) := x"0920";
    tmp(45219) := x"0920";
    tmp(45220) := x"0920";
    tmp(45221) := x"0900";
    tmp(45222) := x"08e0";
    tmp(45223) := x"2141";
    tmp(45224) := x"49a3";
    tmp(45225) := x"61e5";
    tmp(45226) := x"7248";
    tmp(45227) := x"936d";
    tmp(45228) := x"abcf";
    tmp(45229) := x"a3af";
    tmp(45230) := x"a3cf";
    tmp(45231) := x"a3af";
    tmp(45232) := x"abf0";
    tmp(45233) := x"b40f";
    tmp(45234) := x"9b8d";
    tmp(45235) := x"932c";
    tmp(45236) := x"9b4d";
    tmp(45237) := x"9b4d";
    tmp(45238) := x"9b2c";
    tmp(45239) := x"92cb";
    tmp(45240) := x"92aa";
    tmp(45241) := x"9aeb";
    tmp(45242) := x"9b0b";
    tmp(45243) := x"92eb";
    tmp(45244) := x"92cb";
    tmp(45245) := x"92cb";
    tmp(45246) := x"8a6a";
    tmp(45247) := x"7a28";
    tmp(45248) := x"69e6";
    tmp(45249) := x"8a68";
    tmp(45250) := x"8a68";
    tmp(45251) := x"9a88";
    tmp(45252) := x"aac9";
    tmp(45253) := x"aae9";
    tmp(45254) := x"aac9";
    tmp(45255) := x"b309";
    tmp(45256) := x"aae9";
    tmp(45257) := x"bb4b";
    tmp(45258) := x"bb6b";
    tmp(45259) := x"bb4b";
    tmp(45260) := x"b34b";
    tmp(45261) := x"b34b";
    tmp(45262) := x"bb6b";
    tmp(45263) := x"bb8c";
    tmp(45264) := x"c3ae";
    tmp(45265) := x"ab4d";
    tmp(45266) := x"92cb";
    tmp(45267) := x"28c2";
    tmp(45268) := x"1041";
    tmp(45269) := x"28c3";
    tmp(45270) := x"1862";
    tmp(45271) := x"2082";
    tmp(45272) := x"5123";
    tmp(45273) := x"3041";
    tmp(45274) := x"1000";
    tmp(45275) := x"1800";
    tmp(45276) := x"1800";
    tmp(45277) := x"1800";
    tmp(45278) := x"1800";
    tmp(45279) := x"2000";
    tmp(45280) := x"2000";
    tmp(45281) := x"2000";
    tmp(45282) := x"1800";
    tmp(45283) := x"1800";
    tmp(45284) := x"2000";
    tmp(45285) := x"3000";
    tmp(45286) := x"3000";
    tmp(45287) := x"5000";
    tmp(45288) := x"5000";
    tmp(45289) := x"5800";
    tmp(45290) := x"6000";
    tmp(45291) := x"6800";
    tmp(45292) := x"6800";
    tmp(45293) := x"7800";
    tmp(45294) := x"8800";
    tmp(45295) := x"9000";
    tmp(45296) := x"a820";
    tmp(45297) := x"b820";
    tmp(45298) := x"b020";
    tmp(45299) := x"b820";
    tmp(45300) := x"b820";
    tmp(45301) := x"e841";
    tmp(45302) := x"d061";
    tmp(45303) := x"4061";
    tmp(45304) := x"1040";
    tmp(45305) := x"1040";
    tmp(45306) := x"0840";
    tmp(45307) := x"0840";
    tmp(45308) := x"0840";
    tmp(45309) := x"0840";
    tmp(45310) := x"0840";
    tmp(45311) := x"0840";
    tmp(45312) := x"0840";
    tmp(45313) := x"0840";
    tmp(45314) := x"0840";
    tmp(45315) := x"0840";
    tmp(45316) := x"0840";
    tmp(45317) := x"001f";
    tmp(45318) := x"001f";
    tmp(45319) := x"001f";
    tmp(45320) := x"001f";
    tmp(45321) := x"001f";
    tmp(45322) := x"001f";
    tmp(45323) := x"001f";
    tmp(45324) := x"001f";
    tmp(45325) := x"001f";
    tmp(45326) := x"001f";
    tmp(45327) := x"001f";
    tmp(45328) := x"001f";
    tmp(45329) := x"001f";
    tmp(45330) := x"001f";
    tmp(45331) := x"001f";
    tmp(45332) := x"001f";
    tmp(45333) := x"001f";
    tmp(45334) := x"001f";
    tmp(45335) := x"001f";
    tmp(45336) := x"001f";
    tmp(45337) := x"001f";
    tmp(45338) := x"001f";
    tmp(45339) := x"001f";
    tmp(45340) := x"001f";
    tmp(45341) := x"001f";
    tmp(45342) := x"001f";
    tmp(45343) := x"001f";
    tmp(45344) := x"001f";
    tmp(45345) := x"001f";
    tmp(45346) := x"001f";
    tmp(45347) := x"001f";
    tmp(45348) := x"001f";
    tmp(45349) := x"001f";
    tmp(45350) := x"001f";
    tmp(45351) := x"001f";
    tmp(45352) := x"001f";
    tmp(45353) := x"001f";
    tmp(45354) := x"001f";
    tmp(45355) := x"001f";
    tmp(45356) := x"001f";
    tmp(45357) := x"0840";
    tmp(45358) := x"0840";
    tmp(45359) := x"0840";
    tmp(45360) := x"0000";
    tmp(45361) := x"08a0";
    tmp(45362) := x"08a1";
    tmp(45363) := x"08a1";
    tmp(45364) := x"08a1";
    tmp(45365) := x"08a1";
    tmp(45366) := x"08a1";
    tmp(45367) := x"08a1";
    tmp(45368) := x"08a1";
    tmp(45369) := x"08a1";
    tmp(45370) := x"08a1";
    tmp(45371) := x"10a1";
    tmp(45372) := x"10a1";
    tmp(45373) := x"10a1";
    tmp(45374) := x"1081";
    tmp(45375) := x"1081";
    tmp(45376) := x"0881";
    tmp(45377) := x"0881";
    tmp(45378) := x"0881";
    tmp(45379) := x"0860";
    tmp(45380) := x"0860";
    tmp(45381) := x"0860";
    tmp(45382) := x"0860";
    tmp(45383) := x"0860";
    tmp(45384) := x"0860";
    tmp(45385) := x"0860";
    tmp(45386) := x"0860";
    tmp(45387) := x"0860";
    tmp(45388) := x"0860";
    tmp(45389) := x"0860";
    tmp(45390) := x"0860";
    tmp(45391) := x"0860";
    tmp(45392) := x"0860";
    tmp(45393) := x"0860";
    tmp(45394) := x"0860";
    tmp(45395) := x"0860";
    tmp(45396) := x"0860";
    tmp(45397) := x"0860";
    tmp(45398) := x"0860";
    tmp(45399) := x"0860";
    tmp(45400) := x"0860";
    tmp(45401) := x"0860";
    tmp(45402) := x"0860";
    tmp(45403) := x"0880";
    tmp(45404) := x"0880";
    tmp(45405) := x"0880";
    tmp(45406) := x"08a0";
    tmp(45407) := x"08a0";
    tmp(45408) := x"08a0";
    tmp(45409) := x"08c0";
    tmp(45410) := x"08c0";
    tmp(45411) := x"08c0";
    tmp(45412) := x"08c0";
    tmp(45413) := x"08e0";
    tmp(45414) := x"08e0";
    tmp(45415) := x"08e0";
    tmp(45416) := x"08e0";
    tmp(45417) := x"08e0";
    tmp(45418) := x"0900";
    tmp(45419) := x"0900";
    tmp(45420) := x"0920";
    tmp(45421) := x"0920";
    tmp(45422) := x"0920";
    tmp(45423) := x"0920";
    tmp(45424) := x"0920";
    tmp(45425) := x"0920";
    tmp(45426) := x"0920";
    tmp(45427) := x"0900";
    tmp(45428) := x"0920";
    tmp(45429) := x"0900";
    tmp(45430) := x"0900";
    tmp(45431) := x"0900";
    tmp(45432) := x"0900";
    tmp(45433) := x"0900";
    tmp(45434) := x"0900";
    tmp(45435) := x"08e0";
    tmp(45436) := x"08e0";
    tmp(45437) := x"08e0";
    tmp(45438) := x"08e0";
    tmp(45439) := x"08e0";
    tmp(45440) := x"0900";
    tmp(45441) := x"08e0";
    tmp(45442) := x"0900";
    tmp(45443) := x"0900";
    tmp(45444) := x"0900";
    tmp(45445) := x"0900";
    tmp(45446) := x"0900";
    tmp(45447) := x"0900";
    tmp(45448) := x"0900";
    tmp(45449) := x"0900";
    tmp(45450) := x"0920";
    tmp(45451) := x"0920";
    tmp(45452) := x"0920";
    tmp(45453) := x"0920";
    tmp(45454) := x"0920";
    tmp(45455) := x"0920";
    tmp(45456) := x"0920";
    tmp(45457) := x"0920";
    tmp(45458) := x"0920";
    tmp(45459) := x"0920";
    tmp(45460) := x"0920";
    tmp(45461) := x"0900";
    tmp(45462) := x"1100";
    tmp(45463) := x"2942";
    tmp(45464) := x"4184";
    tmp(45465) := x"59e6";
    tmp(45466) := x"7aca";
    tmp(45467) := x"a3cf";
    tmp(45468) := x"938e";
    tmp(45469) := x"938e";
    tmp(45470) := x"936e";
    tmp(45471) := x"8b4d";
    tmp(45472) := x"938e";
    tmp(45473) := x"9bcf";
    tmp(45474) := x"934d";
    tmp(45475) := x"82ec";
    tmp(45476) := x"8b0c";
    tmp(45477) := x"8b0c";
    tmp(45478) := x"8b0c";
    tmp(45479) := x"8aeb";
    tmp(45480) := x"8aaa";
    tmp(45481) := x"8aaa";
    tmp(45482) := x"8acb";
    tmp(45483) := x"7a69";
    tmp(45484) := x"59a6";
    tmp(45485) := x"5186";
    tmp(45486) := x"5186";
    tmp(45487) := x"59a6";
    tmp(45488) := x"61c6";
    tmp(45489) := x"7207";
    tmp(45490) := x"9268";
    tmp(45491) := x"9aa9";
    tmp(45492) := x"a2c9";
    tmp(45493) := x"a2c8";
    tmp(45494) := x"aae9";
    tmp(45495) := x"aaea";
    tmp(45496) := x"a2ca";
    tmp(45497) := x"b34b";
    tmp(45498) := x"bb6c";
    tmp(45499) := x"bb6c";
    tmp(45500) := x"b34b";
    tmp(45501) := x"b36b";
    tmp(45502) := x"b34b";
    tmp(45503) := x"ab2b";
    tmp(45504) := x"b36d";
    tmp(45505) := x"ab6d";
    tmp(45506) := x"82aa";
    tmp(45507) := x"3903";
    tmp(45508) := x"20a2";
    tmp(45509) := x"1882";
    tmp(45510) := x"0841";
    tmp(45511) := x"38e2";
    tmp(45512) := x"3861";
    tmp(45513) := x"1000";
    tmp(45514) := x"1000";
    tmp(45515) := x"1800";
    tmp(45516) := x"2000";
    tmp(45517) := x"1800";
    tmp(45518) := x"2000";
    tmp(45519) := x"3000";
    tmp(45520) := x"2000";
    tmp(45521) := x"2000";
    tmp(45522) := x"2000";
    tmp(45523) := x"2800";
    tmp(45524) := x"3000";
    tmp(45525) := x"3000";
    tmp(45526) := x"3800";
    tmp(45527) := x"4800";
    tmp(45528) := x"5800";
    tmp(45529) := x"5000";
    tmp(45530) := x"6000";
    tmp(45531) := x"6800";
    tmp(45532) := x"7000";
    tmp(45533) := x"7000";
    tmp(45534) := x"8000";
    tmp(45535) := x"8800";
    tmp(45536) := x"9800";
    tmp(45537) := x"a000";
    tmp(45538) := x"b820";
    tmp(45539) := x"b020";
    tmp(45540) := x"a820";
    tmp(45541) := x"d820";
    tmp(45542) := x"f041";
    tmp(45543) := x"8861";
    tmp(45544) := x"1040";
    tmp(45545) := x"1040";
    tmp(45546) := x"1040";
    tmp(45547) := x"0840";
    tmp(45548) := x"0840";
    tmp(45549) := x"0840";
    tmp(45550) := x"0840";
    tmp(45551) := x"0840";
    tmp(45552) := x"0840";
    tmp(45553) := x"0840";
    tmp(45554) := x"0840";
    tmp(45555) := x"0840";
    tmp(45556) := x"0840";
    tmp(45557) := x"001f";
    tmp(45558) := x"001f";
    tmp(45559) := x"001f";
    tmp(45560) := x"001f";
    tmp(45561) := x"001f";
    tmp(45562) := x"001f";
    tmp(45563) := x"001f";
    tmp(45564) := x"001f";
    tmp(45565) := x"001f";
    tmp(45566) := x"001f";
    tmp(45567) := x"001f";
    tmp(45568) := x"001f";
    tmp(45569) := x"001f";
    tmp(45570) := x"001f";
    tmp(45571) := x"001f";
    tmp(45572) := x"001f";
    tmp(45573) := x"001f";
    tmp(45574) := x"001f";
    tmp(45575) := x"001f";
    tmp(45576) := x"001f";
    tmp(45577) := x"001f";
    tmp(45578) := x"001f";
    tmp(45579) := x"001f";
    tmp(45580) := x"001f";
    tmp(45581) := x"001f";
    tmp(45582) := x"001f";
    tmp(45583) := x"001f";
    tmp(45584) := x"001f";
    tmp(45585) := x"001f";
    tmp(45586) := x"001f";
    tmp(45587) := x"001f";
    tmp(45588) := x"001f";
    tmp(45589) := x"001f";
    tmp(45590) := x"001f";
    tmp(45591) := x"001f";
    tmp(45592) := x"001f";
    tmp(45593) := x"001f";
    tmp(45594) := x"001f";
    tmp(45595) := x"001f";
    tmp(45596) := x"001f";
    tmp(45597) := x"0840";
    tmp(45598) := x"0840";
    tmp(45599) := x"0840";
    tmp(45600) := x"0000";
    tmp(45601) := x"08a0";
    tmp(45602) := x"08a1";
    tmp(45603) := x"08a1";
    tmp(45604) := x"08a1";
    tmp(45605) := x"08a1";
    tmp(45606) := x"08a1";
    tmp(45607) := x"08a1";
    tmp(45608) := x"08a1";
    tmp(45609) := x"08a1";
    tmp(45610) := x"08a1";
    tmp(45611) := x"08a1";
    tmp(45612) := x"10a1";
    tmp(45613) := x"10a1";
    tmp(45614) := x"10a1";
    tmp(45615) := x"08a1";
    tmp(45616) := x"08a1";
    tmp(45617) := x"0881";
    tmp(45618) := x"0881";
    tmp(45619) := x"0881";
    tmp(45620) := x"0881";
    tmp(45621) := x"0860";
    tmp(45622) := x"0881";
    tmp(45623) := x"0860";
    tmp(45624) := x"0860";
    tmp(45625) := x"0860";
    tmp(45626) := x"0860";
    tmp(45627) := x"0860";
    tmp(45628) := x"0860";
    tmp(45629) := x"0861";
    tmp(45630) := x"0860";
    tmp(45631) := x"0860";
    tmp(45632) := x"0860";
    tmp(45633) := x"0860";
    tmp(45634) := x"0860";
    tmp(45635) := x"0860";
    tmp(45636) := x"0860";
    tmp(45637) := x"0860";
    tmp(45638) := x"0860";
    tmp(45639) := x"0860";
    tmp(45640) := x"0860";
    tmp(45641) := x"0860";
    tmp(45642) := x"0860";
    tmp(45643) := x"0880";
    tmp(45644) := x"0880";
    tmp(45645) := x"0880";
    tmp(45646) := x"0880";
    tmp(45647) := x"08a0";
    tmp(45648) := x"08a0";
    tmp(45649) := x"08a0";
    tmp(45650) := x"08a0";
    tmp(45651) := x"08c0";
    tmp(45652) := x"08c0";
    tmp(45653) := x"08c0";
    tmp(45654) := x"08e0";
    tmp(45655) := x"08e0";
    tmp(45656) := x"08e0";
    tmp(45657) := x"08e0";
    tmp(45658) := x"08e0";
    tmp(45659) := x"0900";
    tmp(45660) := x"0900";
    tmp(45661) := x"0920";
    tmp(45662) := x"0920";
    tmp(45663) := x"0900";
    tmp(45664) := x"0920";
    tmp(45665) := x"0920";
    tmp(45666) := x"0920";
    tmp(45667) := x"0920";
    tmp(45668) := x"0900";
    tmp(45669) := x"0900";
    tmp(45670) := x"0900";
    tmp(45671) := x"0900";
    tmp(45672) := x"0900";
    tmp(45673) := x"0900";
    tmp(45674) := x"0900";
    tmp(45675) := x"0900";
    tmp(45676) := x"08e0";
    tmp(45677) := x"08e0";
    tmp(45678) := x"08e0";
    tmp(45679) := x"08e0";
    tmp(45680) := x"08e0";
    tmp(45681) := x"08e0";
    tmp(45682) := x"0900";
    tmp(45683) := x"0900";
    tmp(45684) := x"0900";
    tmp(45685) := x"0900";
    tmp(45686) := x"0900";
    tmp(45687) := x"0900";
    tmp(45688) := x"0900";
    tmp(45689) := x"0920";
    tmp(45690) := x"0920";
    tmp(45691) := x"0920";
    tmp(45692) := x"0920";
    tmp(45693) := x"0920";
    tmp(45694) := x"0920";
    tmp(45695) := x"0920";
    tmp(45696) := x"0920";
    tmp(45697) := x"0920";
    tmp(45698) := x"0940";
    tmp(45699) := x"0920";
    tmp(45700) := x"0920";
    tmp(45701) := x"0900";
    tmp(45702) := x"18e1";
    tmp(45703) := x"2102";
    tmp(45704) := x"3964";
    tmp(45705) := x"49c6";
    tmp(45706) := x"8b4d";
    tmp(45707) := x"936e";
    tmp(45708) := x"8b4d";
    tmp(45709) := x"7b0c";
    tmp(45710) := x"72cb";
    tmp(45711) := x"72cb";
    tmp(45712) := x"7aec";
    tmp(45713) := x"7aec";
    tmp(45714) := x"72cb";
    tmp(45715) := x"6a8a";
    tmp(45716) := x"6a69";
    tmp(45717) := x"6a8a";
    tmp(45718) := x"72a9";
    tmp(45719) := x"6a69";
    tmp(45720) := x"6a48";
    tmp(45721) := x"59c6";
    tmp(45722) := x"5185";
    tmp(45723) := x"3924";
    tmp(45724) := x"4124";
    tmp(45725) := x"5186";
    tmp(45726) := x"6a08";
    tmp(45727) := x"7a49";
    tmp(45728) := x"7a48";
    tmp(45729) := x"8268";
    tmp(45730) := x"92ca";
    tmp(45731) := x"92a9";
    tmp(45732) := x"9288";
    tmp(45733) := x"9aa9";
    tmp(45734) := x"9aa9";
    tmp(45735) := x"aaea";
    tmp(45736) := x"ab2a";
    tmp(45737) := x"9ac9";
    tmp(45738) := x"ab4a";
    tmp(45739) := x"b34b";
    tmp(45740) := x"ab2b";
    tmp(45741) := x"ab4a";
    tmp(45742) := x"a34b";
    tmp(45743) := x"9b2b";
    tmp(45744) := x"92eb";
    tmp(45745) := x"828a";
    tmp(45746) := x"4965";
    tmp(45747) := x"20a2";
    tmp(45748) := x"1041";
    tmp(45749) := x"0820";
    tmp(45750) := x"0841";
    tmp(45751) := x"3081";
    tmp(45752) := x"2020";
    tmp(45753) := x"1000";
    tmp(45754) := x"1000";
    tmp(45755) := x"1800";
    tmp(45756) := x"1800";
    tmp(45757) := x"1800";
    tmp(45758) := x"2000";
    tmp(45759) := x"2000";
    tmp(45760) := x"2000";
    tmp(45761) := x"2000";
    tmp(45762) := x"1800";
    tmp(45763) := x"2000";
    tmp(45764) := x"2800";
    tmp(45765) := x"3000";
    tmp(45766) := x"3800";
    tmp(45767) := x"4000";
    tmp(45768) := x"5000";
    tmp(45769) := x"5800";
    tmp(45770) := x"6000";
    tmp(45771) := x"7000";
    tmp(45772) := x"8800";
    tmp(45773) := x"8000";
    tmp(45774) := x"9020";
    tmp(45775) := x"9820";
    tmp(45776) := x"8800";
    tmp(45777) := x"9800";
    tmp(45778) := x"b020";
    tmp(45779) := x"b020";
    tmp(45780) := x"a800";
    tmp(45781) := x"b020";
    tmp(45782) := x"d820";
    tmp(45783) := x"c861";
    tmp(45784) := x"3040";
    tmp(45785) := x"1040";
    tmp(45786) := x"0840";
    tmp(45787) := x"0840";
    tmp(45788) := x"0840";
    tmp(45789) := x"0840";
    tmp(45790) := x"0840";
    tmp(45791) := x"0840";
    tmp(45792) := x"0840";
    tmp(45793) := x"0840";
    tmp(45794) := x"0840";
    tmp(45795) := x"0840";
    tmp(45796) := x"0840";
    tmp(45797) := x"001f";
    tmp(45798) := x"001f";
    tmp(45799) := x"001f";
    tmp(45800) := x"001f";
    tmp(45801) := x"001f";
    tmp(45802) := x"001f";
    tmp(45803) := x"001f";
    tmp(45804) := x"001f";
    tmp(45805) := x"001f";
    tmp(45806) := x"001f";
    tmp(45807) := x"001f";
    tmp(45808) := x"001f";
    tmp(45809) := x"001f";
    tmp(45810) := x"001f";
    tmp(45811) := x"001f";
    tmp(45812) := x"001f";
    tmp(45813) := x"001f";
    tmp(45814) := x"001f";
    tmp(45815) := x"001f";
    tmp(45816) := x"001f";
    tmp(45817) := x"001f";
    tmp(45818) := x"001f";
    tmp(45819) := x"001f";
    tmp(45820) := x"001f";
    tmp(45821) := x"001f";
    tmp(45822) := x"001f";
    tmp(45823) := x"001f";
    tmp(45824) := x"001f";
    tmp(45825) := x"001f";
    tmp(45826) := x"001f";
    tmp(45827) := x"001f";
    tmp(45828) := x"001f";
    tmp(45829) := x"001f";
    tmp(45830) := x"001f";
    tmp(45831) := x"001f";
    tmp(45832) := x"001f";
    tmp(45833) := x"001f";
    tmp(45834) := x"001f";
    tmp(45835) := x"001f";
    tmp(45836) := x"001f";
    tmp(45837) := x"0840";
    tmp(45838) := x"0840";
    tmp(45839) := x"0840";
    tmp(45840) := x"0000";
    tmp(45841) := x"08a0";
    tmp(45842) := x"08a0";
    tmp(45843) := x"08c1";
    tmp(45844) := x"08c1";
    tmp(45845) := x"08a1";
    tmp(45846) := x"08c1";
    tmp(45847) := x"08a1";
    tmp(45848) := x"08a1";
    tmp(45849) := x"08a1";
    tmp(45850) := x"10a1";
    tmp(45851) := x"08a1";
    tmp(45852) := x"10a1";
    tmp(45853) := x"08a1";
    tmp(45854) := x"10a1";
    tmp(45855) := x"10a1";
    tmp(45856) := x"10a1";
    tmp(45857) := x"08a1";
    tmp(45858) := x"08a1";
    tmp(45859) := x"0881";
    tmp(45860) := x"0881";
    tmp(45861) := x"0881";
    tmp(45862) := x"0881";
    tmp(45863) := x"0880";
    tmp(45864) := x"0860";
    tmp(45865) := x"0860";
    tmp(45866) := x"0881";
    tmp(45867) := x"0861";
    tmp(45868) := x"0860";
    tmp(45869) := x"1081";
    tmp(45870) := x"1061";
    tmp(45871) := x"1061";
    tmp(45872) := x"0861";
    tmp(45873) := x"0861";
    tmp(45874) := x"0860";
    tmp(45875) := x"0860";
    tmp(45876) := x"0860";
    tmp(45877) := x"0860";
    tmp(45878) := x"0860";
    tmp(45879) := x"0860";
    tmp(45880) := x"0860";
    tmp(45881) := x"0860";
    tmp(45882) := x"0860";
    tmp(45883) := x"0860";
    tmp(45884) := x"0880";
    tmp(45885) := x"0880";
    tmp(45886) := x"0880";
    tmp(45887) := x"0880";
    tmp(45888) := x"08a0";
    tmp(45889) := x"08a0";
    tmp(45890) := x"08a0";
    tmp(45891) := x"08a0";
    tmp(45892) := x"08c0";
    tmp(45893) := x"08c0";
    tmp(45894) := x"08c0";
    tmp(45895) := x"08c0";
    tmp(45896) := x"08c0";
    tmp(45897) := x"08e0";
    tmp(45898) := x"08e0";
    tmp(45899) := x"08e0";
    tmp(45900) := x"0900";
    tmp(45901) := x"0900";
    tmp(45902) := x"0900";
    tmp(45903) := x"0900";
    tmp(45904) := x"0900";
    tmp(45905) := x"0900";
    tmp(45906) := x"0900";
    tmp(45907) := x"0920";
    tmp(45908) := x"0900";
    tmp(45909) := x"0900";
    tmp(45910) := x"0900";
    tmp(45911) := x"0900";
    tmp(45912) := x"0900";
    tmp(45913) := x"0900";
    tmp(45914) := x"0900";
    tmp(45915) := x"0900";
    tmp(45916) := x"08e0";
    tmp(45917) := x"08e0";
    tmp(45918) := x"08e0";
    tmp(45919) := x"08e0";
    tmp(45920) := x"08e0";
    tmp(45921) := x"08e0";
    tmp(45922) := x"08e0";
    tmp(45923) := x"08e0";
    tmp(45924) := x"0900";
    tmp(45925) := x"0900";
    tmp(45926) := x"0900";
    tmp(45927) := x"0900";
    tmp(45928) := x"0900";
    tmp(45929) := x"0920";
    tmp(45930) := x"0900";
    tmp(45931) := x"0920";
    tmp(45932) := x"0920";
    tmp(45933) := x"0920";
    tmp(45934) := x"0920";
    tmp(45935) := x"0920";
    tmp(45936) := x"0920";
    tmp(45937) := x"0920";
    tmp(45938) := x"0920";
    tmp(45939) := x"0920";
    tmp(45940) := x"0920";
    tmp(45941) := x"10a0";
    tmp(45942) := x"1081";
    tmp(45943) := x"18a2";
    tmp(45944) := x"2924";
    tmp(45945) := x"41a6";
    tmp(45946) := x"730c";
    tmp(45947) := x"730c";
    tmp(45948) := x"628a";
    tmp(45949) := x"5a49";
    tmp(45950) := x"5228";
    tmp(45951) := x"5208";
    tmp(45952) := x"4a08";
    tmp(45953) := x"41e7";
    tmp(45954) := x"41a6";
    tmp(45955) := x"3165";
    tmp(45956) := x"3144";
    tmp(45957) := x"2904";
    tmp(45958) := x"2924";
    tmp(45959) := x"3124";
    tmp(45960) := x"28c2";
    tmp(45961) := x"1861";
    tmp(45962) := x"30e3";
    tmp(45963) := x"51a6";
    tmp(45964) := x"5a07";
    tmp(45965) := x"6a29";
    tmp(45966) := x"7269";
    tmp(45967) := x"7a69";
    tmp(45968) := x"7228";
    tmp(45969) := x"7248";
    tmp(45970) := x"7a69";
    tmp(45971) := x"8289";
    tmp(45972) := x"8a88";
    tmp(45973) := x"8aa9";
    tmp(45974) := x"92c9";
    tmp(45975) := x"9aea";
    tmp(45976) := x"92ea";
    tmp(45977) := x"92e9";
    tmp(45978) := x"92c9";
    tmp(45979) := x"92ca";
    tmp(45980) := x"92c9";
    tmp(45981) := x"92c9";
    tmp(45982) := x"8ac9";
    tmp(45983) := x"82a9";
    tmp(45984) := x"7a68";
    tmp(45985) := x"3924";
    tmp(45986) := x"1041";
    tmp(45987) := x"0000";
    tmp(45988) := x"0000";
    tmp(45989) := x"0000";
    tmp(45990) := x"1041";
    tmp(45991) := x"40a2";
    tmp(45992) := x"1000";
    tmp(45993) := x"1000";
    tmp(45994) := x"1000";
    tmp(45995) := x"1000";
    tmp(45996) := x"1800";
    tmp(45997) := x"1800";
    tmp(45998) := x"1800";
    tmp(45999) := x"2000";
    tmp(46000) := x"2800";
    tmp(46001) := x"2000";
    tmp(46002) := x"2000";
    tmp(46003) := x"2000";
    tmp(46004) := x"2800";
    tmp(46005) := x"3000";
    tmp(46006) := x"3000";
    tmp(46007) := x"4000";
    tmp(46008) := x"5000";
    tmp(46009) := x"6000";
    tmp(46010) := x"6800";
    tmp(46011) := x"7800";
    tmp(46012) := x"9020";
    tmp(46013) := x"9020";
    tmp(46014) := x"9020";
    tmp(46015) := x"9020";
    tmp(46016) := x"b020";
    tmp(46017) := x"a000";
    tmp(46018) := x"b800";
    tmp(46019) := x"b020";
    tmp(46020) := x"a820";
    tmp(46021) := x"b820";
    tmp(46022) := x"c020";
    tmp(46023) := x"d041";
    tmp(46024) := x"6861";
    tmp(46025) := x"1840";
    tmp(46026) := x"1040";
    tmp(46027) := x"0840";
    tmp(46028) := x"0840";
    tmp(46029) := x"0840";
    tmp(46030) := x"0840";
    tmp(46031) := x"0840";
    tmp(46032) := x"0840";
    tmp(46033) := x"0840";
    tmp(46034) := x"0840";
    tmp(46035) := x"0840";
    tmp(46036) := x"0840";
    tmp(46037) := x"001f";
    tmp(46038) := x"001f";
    tmp(46039) := x"001f";
    tmp(46040) := x"001f";
    tmp(46041) := x"001f";
    tmp(46042) := x"001f";
    tmp(46043) := x"001f";
    tmp(46044) := x"001f";
    tmp(46045) := x"001f";
    tmp(46046) := x"001f";
    tmp(46047) := x"001f";
    tmp(46048) := x"001f";
    tmp(46049) := x"001f";
    tmp(46050) := x"001f";
    tmp(46051) := x"001f";
    tmp(46052) := x"001f";
    tmp(46053) := x"001f";
    tmp(46054) := x"001f";
    tmp(46055) := x"001f";
    tmp(46056) := x"001f";
    tmp(46057) := x"001f";
    tmp(46058) := x"001f";
    tmp(46059) := x"001f";
    tmp(46060) := x"001f";
    tmp(46061) := x"001f";
    tmp(46062) := x"001f";
    tmp(46063) := x"001f";
    tmp(46064) := x"001f";
    tmp(46065) := x"001f";
    tmp(46066) := x"001f";
    tmp(46067) := x"001f";
    tmp(46068) := x"001f";
    tmp(46069) := x"001f";
    tmp(46070) := x"001f";
    tmp(46071) := x"001f";
    tmp(46072) := x"001f";
    tmp(46073) := x"001f";
    tmp(46074) := x"001f";
    tmp(46075) := x"001f";
    tmp(46076) := x"001f";
    tmp(46077) := x"0840";
    tmp(46078) := x"0840";
    tmp(46079) := x"0840";
    tmp(46080) := x"0000";
    tmp(46081) := x"08c0";
    tmp(46082) := x"08a0";
    tmp(46083) := x"08a1";
    tmp(46084) := x"08c1";
    tmp(46085) := x"08c1";
    tmp(46086) := x"08c1";
    tmp(46087) := x"08c1";
    tmp(46088) := x"10c1";
    tmp(46089) := x"10c1";
    tmp(46090) := x"08c1";
    tmp(46091) := x"10c1";
    tmp(46092) := x"10c1";
    tmp(46093) := x"10a1";
    tmp(46094) := x"10a1";
    tmp(46095) := x"10a1";
    tmp(46096) := x"10a1";
    tmp(46097) := x"10a1";
    tmp(46098) := x"10a1";
    tmp(46099) := x"10a1";
    tmp(46100) := x"08a1";
    tmp(46101) := x"0881";
    tmp(46102) := x"0881";
    tmp(46103) := x"0881";
    tmp(46104) := x"0881";
    tmp(46105) := x"0881";
    tmp(46106) := x"0881";
    tmp(46107) := x"1081";
    tmp(46108) := x"1081";
    tmp(46109) := x"1081";
    tmp(46110) := x"1081";
    tmp(46111) := x"1081";
    tmp(46112) := x"1081";
    tmp(46113) := x"1081";
    tmp(46114) := x"1061";
    tmp(46115) := x"0861";
    tmp(46116) := x"0861";
    tmp(46117) := x"0860";
    tmp(46118) := x"0860";
    tmp(46119) := x"0860";
    tmp(46120) := x"0860";
    tmp(46121) := x"0860";
    tmp(46122) := x"0860";
    tmp(46123) := x"0860";
    tmp(46124) := x"0860";
    tmp(46125) := x"0860";
    tmp(46126) := x"0880";
    tmp(46127) := x"0880";
    tmp(46128) := x"0880";
    tmp(46129) := x"08a0";
    tmp(46130) := x"08a0";
    tmp(46131) := x"08a0";
    tmp(46132) := x"08a0";
    tmp(46133) := x"08c0";
    tmp(46134) := x"08c0";
    tmp(46135) := x"08c0";
    tmp(46136) := x"08c0";
    tmp(46137) := x"08e0";
    tmp(46138) := x"08e0";
    tmp(46139) := x"08e0";
    tmp(46140) := x"08e0";
    tmp(46141) := x"0900";
    tmp(46142) := x"0900";
    tmp(46143) := x"0900";
    tmp(46144) := x"0900";
    tmp(46145) := x"0900";
    tmp(46146) := x"0900";
    tmp(46147) := x"0900";
    tmp(46148) := x"0900";
    tmp(46149) := x"0900";
    tmp(46150) := x"0900";
    tmp(46151) := x"0900";
    tmp(46152) := x"08e0";
    tmp(46153) := x"08e0";
    tmp(46154) := x"0900";
    tmp(46155) := x"08e0";
    tmp(46156) := x"08e0";
    tmp(46157) := x"08e0";
    tmp(46158) := x"08e0";
    tmp(46159) := x"08e0";
    tmp(46160) := x"08e0";
    tmp(46161) := x"08e0";
    tmp(46162) := x"08e0";
    tmp(46163) := x"0900";
    tmp(46164) := x"0900";
    tmp(46165) := x"08e0";
    tmp(46166) := x"0900";
    tmp(46167) := x"0900";
    tmp(46168) := x"0900";
    tmp(46169) := x"0900";
    tmp(46170) := x"0900";
    tmp(46171) := x"0900";
    tmp(46172) := x"0920";
    tmp(46173) := x"0920";
    tmp(46174) := x"0900";
    tmp(46175) := x"0900";
    tmp(46176) := x"0920";
    tmp(46177) := x"0920";
    tmp(46178) := x"0920";
    tmp(46179) := x"0920";
    tmp(46180) := x"08e0";
    tmp(46181) := x"0861";
    tmp(46182) := x"0841";
    tmp(46183) := x"1062";
    tmp(46184) := x"18c3";
    tmp(46185) := x"4a07";
    tmp(46186) := x"4a08";
    tmp(46187) := x"41c7";
    tmp(46188) := x"3185";
    tmp(46189) := x"2945";
    tmp(46190) := x"2945";
    tmp(46191) := x"3186";
    tmp(46192) := x"2945";
    tmp(46193) := x"18a3";
    tmp(46194) := x"1082";
    tmp(46195) := x"1082";
    tmp(46196) := x"1061";
    tmp(46197) := x"1061";
    tmp(46198) := x"1061";
    tmp(46199) := x"1061";
    tmp(46200) := x"1061";
    tmp(46201) := x"20c2";
    tmp(46202) := x"3144";
    tmp(46203) := x"49c7";
    tmp(46204) := x"5a29";
    tmp(46205) := x"6229";
    tmp(46206) := x"6229";
    tmp(46207) := x"5a08";
    tmp(46208) := x"51e7";
    tmp(46209) := x"59e7";
    tmp(46210) := x"6227";
    tmp(46211) := x"7269";
    tmp(46212) := x"7a69";
    tmp(46213) := x"7a68";
    tmp(46214) := x"7a69";
    tmp(46215) := x"7a89";
    tmp(46216) := x"8289";
    tmp(46217) := x"8289";
    tmp(46218) := x"8aea";
    tmp(46219) := x"7248";
    tmp(46220) := x"6207";
    tmp(46221) := x"5185";
    tmp(46222) := x"4144";
    tmp(46223) := x"3924";
    tmp(46224) := x"20a2";
    tmp(46225) := x"1041";
    tmp(46226) := x"0820";
    tmp(46227) := x"0020";
    tmp(46228) := x"0000";
    tmp(46229) := x"0000";
    tmp(46230) := x"5164";
    tmp(46231) := x"3061";
    tmp(46232) := x"1800";
    tmp(46233) := x"1000";
    tmp(46234) := x"1800";
    tmp(46235) := x"1800";
    tmp(46236) := x"2000";
    tmp(46237) := x"1800";
    tmp(46238) := x"1800";
    tmp(46239) := x"2000";
    tmp(46240) := x"2000";
    tmp(46241) := x"2000";
    tmp(46242) := x"2000";
    tmp(46243) := x"2000";
    tmp(46244) := x"2800";
    tmp(46245) := x"2800";
    tmp(46246) := x"3000";
    tmp(46247) := x"3800";
    tmp(46248) := x"5000";
    tmp(46249) := x"5000";
    tmp(46250) := x"6000";
    tmp(46251) := x"7000";
    tmp(46252) := x"8820";
    tmp(46253) := x"9020";
    tmp(46254) := x"8820";
    tmp(46255) := x"8820";
    tmp(46256) := x"a820";
    tmp(46257) := x"b820";
    tmp(46258) := x"a800";
    tmp(46259) := x"a820";
    tmp(46260) := x"a820";
    tmp(46261) := x"b820";
    tmp(46262) := x"b820";
    tmp(46263) := x"f841";
    tmp(46264) := x"b861";
    tmp(46265) := x"3840";
    tmp(46266) := x"1040";
    tmp(46267) := x"0840";
    tmp(46268) := x"0840";
    tmp(46269) := x"0840";
    tmp(46270) := x"0840";
    tmp(46271) := x"0840";
    tmp(46272) := x"0840";
    tmp(46273) := x"0840";
    tmp(46274) := x"0840";
    tmp(46275) := x"0840";
    tmp(46276) := x"0840";
    tmp(46277) := x"001f";
    tmp(46278) := x"001f";
    tmp(46279) := x"001f";
    tmp(46280) := x"001f";
    tmp(46281) := x"001f";
    tmp(46282) := x"001f";
    tmp(46283) := x"001f";
    tmp(46284) := x"001f";
    tmp(46285) := x"001f";
    tmp(46286) := x"001f";
    tmp(46287) := x"001f";
    tmp(46288) := x"001f";
    tmp(46289) := x"001f";
    tmp(46290) := x"001f";
    tmp(46291) := x"001f";
    tmp(46292) := x"001f";
    tmp(46293) := x"001f";
    tmp(46294) := x"001f";
    tmp(46295) := x"001f";
    tmp(46296) := x"001f";
    tmp(46297) := x"001f";
    tmp(46298) := x"001f";
    tmp(46299) := x"001f";
    tmp(46300) := x"001f";
    tmp(46301) := x"001f";
    tmp(46302) := x"001f";
    tmp(46303) := x"001f";
    tmp(46304) := x"001f";
    tmp(46305) := x"001f";
    tmp(46306) := x"001f";
    tmp(46307) := x"001f";
    tmp(46308) := x"001f";
    tmp(46309) := x"001f";
    tmp(46310) := x"001f";
    tmp(46311) := x"001f";
    tmp(46312) := x"001f";
    tmp(46313) := x"001f";
    tmp(46314) := x"001f";
    tmp(46315) := x"001f";
    tmp(46316) := x"001f";
    tmp(46317) := x"0840";
    tmp(46318) := x"1040";
    tmp(46319) := x"0840";
    tmp(46320) := x"0020";
    tmp(46321) := x"08c0";
    tmp(46322) := x"08c0";
    tmp(46323) := x"08a0";
    tmp(46324) := x"08c1";
    tmp(46325) := x"08c1";
    tmp(46326) := x"08e1";
    tmp(46327) := x"08e1";
    tmp(46328) := x"10e1";
    tmp(46329) := x"10e1";
    tmp(46330) := x"10c1";
    tmp(46331) := x"10c1";
    tmp(46332) := x"10c1";
    tmp(46333) := x"10c1";
    tmp(46334) := x"10c1";
    tmp(46335) := x"10c1";
    tmp(46336) := x"10c1";
    tmp(46337) := x"10a1";
    tmp(46338) := x"10a1";
    tmp(46339) := x"10a1";
    tmp(46340) := x"10a1";
    tmp(46341) := x"10a1";
    tmp(46342) := x"08a1";
    tmp(46343) := x"08a1";
    tmp(46344) := x"0881";
    tmp(46345) := x"0881";
    tmp(46346) := x"0881";
    tmp(46347) := x"0881";
    tmp(46348) := x"1081";
    tmp(46349) := x"1081";
    tmp(46350) := x"1081";
    tmp(46351) := x"1081";
    tmp(46352) := x"1081";
    tmp(46353) := x"1081";
    tmp(46354) := x"1081";
    tmp(46355) := x"1081";
    tmp(46356) := x"0861";
    tmp(46357) := x"0861";
    tmp(46358) := x"0860";
    tmp(46359) := x"0860";
    tmp(46360) := x"0860";
    tmp(46361) := x"0860";
    tmp(46362) := x"0860";
    tmp(46363) := x"0860";
    tmp(46364) := x"0860";
    tmp(46365) := x"0860";
    tmp(46366) := x"0860";
    tmp(46367) := x"0880";
    tmp(46368) := x"0880";
    tmp(46369) := x"0880";
    tmp(46370) := x"08a0";
    tmp(46371) := x"08a0";
    tmp(46372) := x"08a0";
    tmp(46373) := x"08a0";
    tmp(46374) := x"08c0";
    tmp(46375) := x"08c0";
    tmp(46376) := x"08c0";
    tmp(46377) := x"08c0";
    tmp(46378) := x"08e0";
    tmp(46379) := x"08c0";
    tmp(46380) := x"08e0";
    tmp(46381) := x"08e0";
    tmp(46382) := x"08e0";
    tmp(46383) := x"08e0";
    tmp(46384) := x"08e0";
    tmp(46385) := x"0900";
    tmp(46386) := x"0900";
    tmp(46387) := x"0900";
    tmp(46388) := x"0900";
    tmp(46389) := x"0900";
    tmp(46390) := x"08e0";
    tmp(46391) := x"08e0";
    tmp(46392) := x"08e0";
    tmp(46393) := x"08e0";
    tmp(46394) := x"08e0";
    tmp(46395) := x"08c0";
    tmp(46396) := x"08e0";
    tmp(46397) := x"08e0";
    tmp(46398) := x"08e0";
    tmp(46399) := x"08e0";
    tmp(46400) := x"08e0";
    tmp(46401) := x"08e0";
    tmp(46402) := x"08e0";
    tmp(46403) := x"08e0";
    tmp(46404) := x"08e0";
    tmp(46405) := x"08e0";
    tmp(46406) := x"0900";
    tmp(46407) := x"0900";
    tmp(46408) := x"0900";
    tmp(46409) := x"0900";
    tmp(46410) := x"0900";
    tmp(46411) := x"0900";
    tmp(46412) := x"0900";
    tmp(46413) := x"0900";
    tmp(46414) := x"0920";
    tmp(46415) := x"0900";
    tmp(46416) := x"0920";
    tmp(46417) := x"0920";
    tmp(46418) := x"0920";
    tmp(46419) := x"0900";
    tmp(46420) := x"0880";
    tmp(46421) := x"0841";
    tmp(46422) := x"0841";
    tmp(46423) := x"0861";
    tmp(46424) := x"18e3";
    tmp(46425) := x"2104";
    tmp(46426) := x"2104";
    tmp(46427) := x"18a3";
    tmp(46428) := x"10a2";
    tmp(46429) := x"1082";
    tmp(46430) := x"10a2";
    tmp(46431) := x"2104";
    tmp(46432) := x"18a2";
    tmp(46433) := x"1061";
    tmp(46434) := x"0841";
    tmp(46435) := x"0841";
    tmp(46436) := x"0821";
    tmp(46437) := x"0821";
    tmp(46438) := x"0841";
    tmp(46439) := x"0861";
    tmp(46440) := x"10a2";
    tmp(46441) := x"18c3";
    tmp(46442) := x"18c3";
    tmp(46443) := x"2104";
    tmp(46444) := x"3145";
    tmp(46445) := x"3166";
    tmp(46446) := x"2925";
    tmp(46447) := x"20e4";
    tmp(46448) := x"20e4";
    tmp(46449) := x"2104";
    tmp(46450) := x"2924";
    tmp(46451) := x"3965";
    tmp(46452) := x"3965";
    tmp(46453) := x"3965";
    tmp(46454) := x"3965";
    tmp(46455) := x"3965";
    tmp(46456) := x"3124";
    tmp(46457) := x"28e3";
    tmp(46458) := x"20a2";
    tmp(46459) := x"20a2";
    tmp(46460) := x"1861";
    tmp(46461) := x"1041";
    tmp(46462) := x"0820";
    tmp(46463) := x"0820";
    tmp(46464) := x"0820";
    tmp(46465) := x"0820";
    tmp(46466) := x"0000";
    tmp(46467) := x"0020";
    tmp(46468) := x"0000";
    tmp(46469) := x"0820";
    tmp(46470) := x"5944";
    tmp(46471) := x"2020";
    tmp(46472) := x"1800";
    tmp(46473) := x"1800";
    tmp(46474) := x"1000";
    tmp(46475) := x"1800";
    tmp(46476) := x"2000";
    tmp(46477) := x"2000";
    tmp(46478) := x"2000";
    tmp(46479) := x"2800";
    tmp(46480) := x"5861";
    tmp(46481) := x"5061";
    tmp(46482) := x"2000";
    tmp(46483) := x"2000";
    tmp(46484) := x"2000";
    tmp(46485) := x"2800";
    tmp(46486) := x"3000";
    tmp(46487) := x"3800";
    tmp(46488) := x"4000";
    tmp(46489) := x"5000";
    tmp(46490) := x"6000";
    tmp(46491) := x"7000";
    tmp(46492) := x"8000";
    tmp(46493) := x"8800";
    tmp(46494) := x"8800";
    tmp(46495) := x"8800";
    tmp(46496) := x"a020";
    tmp(46497) := x"b020";
    tmp(46498) := x"a800";
    tmp(46499) := x"b020";
    tmp(46500) := x"b820";
    tmp(46501) := x"b820";
    tmp(46502) := x"c820";
    tmp(46503) := x"e041";
    tmp(46504) := x"f061";
    tmp(46505) := x"8861";
    tmp(46506) := x"1840";
    tmp(46507) := x"1040";
    tmp(46508) := x"1040";
    tmp(46509) := x"0840";
    tmp(46510) := x"0840";
    tmp(46511) := x"0840";
    tmp(46512) := x"0840";
    tmp(46513) := x"0840";
    tmp(46514) := x"0840";
    tmp(46515) := x"0840";
    tmp(46516) := x"0840";
    tmp(46517) := x"001f";
    tmp(46518) := x"001f";
    tmp(46519) := x"001f";
    tmp(46520) := x"001f";
    tmp(46521) := x"001f";
    tmp(46522) := x"001f";
    tmp(46523) := x"001f";
    tmp(46524) := x"001f";
    tmp(46525) := x"001f";
    tmp(46526) := x"001f";
    tmp(46527) := x"001f";
    tmp(46528) := x"001f";
    tmp(46529) := x"001f";
    tmp(46530) := x"001f";
    tmp(46531) := x"001f";
    tmp(46532) := x"001f";
    tmp(46533) := x"001f";
    tmp(46534) := x"001f";
    tmp(46535) := x"001f";
    tmp(46536) := x"001f";
    tmp(46537) := x"001f";
    tmp(46538) := x"001f";
    tmp(46539) := x"001f";
    tmp(46540) := x"001f";
    tmp(46541) := x"001f";
    tmp(46542) := x"001f";
    tmp(46543) := x"001f";
    tmp(46544) := x"001f";
    tmp(46545) := x"001f";
    tmp(46546) := x"001f";
    tmp(46547) := x"001f";
    tmp(46548) := x"001f";
    tmp(46549) := x"001f";
    tmp(46550) := x"001f";
    tmp(46551) := x"001f";
    tmp(46552) := x"001f";
    tmp(46553) := x"001f";
    tmp(46554) := x"001f";
    tmp(46555) := x"001f";
    tmp(46556) := x"001f";
    tmp(46557) := x"1040";
    tmp(46558) := x"0840";
    tmp(46559) := x"0840";
    tmp(46560) := x"0020";
    tmp(46561) := x"08c0";
    tmp(46562) := x"08c0";
    tmp(46563) := x"08c0";
    tmp(46564) := x"08c1";
    tmp(46565) := x"08c1";
    tmp(46566) := x"08e1";
    tmp(46567) := x"10e1";
    tmp(46568) := x"10e1";
    tmp(46569) := x"1101";
    tmp(46570) := x"10e1";
    tmp(46571) := x"10e1";
    tmp(46572) := x"10e1";
    tmp(46573) := x"10c1";
    tmp(46574) := x"10e1";
    tmp(46575) := x"10c1";
    tmp(46576) := x"10c1";
    tmp(46577) := x"10c1";
    tmp(46578) := x"10c1";
    tmp(46579) := x"10a1";
    tmp(46580) := x"10a1";
    tmp(46581) := x"10a1";
    tmp(46582) := x"10a1";
    tmp(46583) := x"08a1";
    tmp(46584) := x"0881";
    tmp(46585) := x"0881";
    tmp(46586) := x"0881";
    tmp(46587) := x"1081";
    tmp(46588) := x"1081";
    tmp(46589) := x"1081";
    tmp(46590) := x"1081";
    tmp(46591) := x"1081";
    tmp(46592) := x"1081";
    tmp(46593) := x"1081";
    tmp(46594) := x"1081";
    tmp(46595) := x"1081";
    tmp(46596) := x"1061";
    tmp(46597) := x"0861";
    tmp(46598) := x"0861";
    tmp(46599) := x"0861";
    tmp(46600) := x"0860";
    tmp(46601) := x"0860";
    tmp(46602) := x"0860";
    tmp(46603) := x"0860";
    tmp(46604) := x"0860";
    tmp(46605) := x"0860";
    tmp(46606) := x"0860";
    tmp(46607) := x"0860";
    tmp(46608) := x"0880";
    tmp(46609) := x"0880";
    tmp(46610) := x"0880";
    tmp(46611) := x"08a0";
    tmp(46612) := x"08a0";
    tmp(46613) := x"08a0";
    tmp(46614) := x"08a0";
    tmp(46615) := x"08a0";
    tmp(46616) := x"08c0";
    tmp(46617) := x"08c0";
    tmp(46618) := x"08c0";
    tmp(46619) := x"08c0";
    tmp(46620) := x"08c0";
    tmp(46621) := x"08e0";
    tmp(46622) := x"08e0";
    tmp(46623) := x"08e0";
    tmp(46624) := x"08e0";
    tmp(46625) := x"08e0";
    tmp(46626) := x"08e0";
    tmp(46627) := x"08e0";
    tmp(46628) := x"08e0";
    tmp(46629) := x"08e0";
    tmp(46630) := x"08e0";
    tmp(46631) := x"08e0";
    tmp(46632) := x"08e0";
    tmp(46633) := x"08c0";
    tmp(46634) := x"08e0";
    tmp(46635) := x"08c0";
    tmp(46636) := x"08c0";
    tmp(46637) := x"08e0";
    tmp(46638) := x"08e0";
    tmp(46639) := x"08e0";
    tmp(46640) := x"08e0";
    tmp(46641) := x"08e0";
    tmp(46642) := x"08e0";
    tmp(46643) := x"08e0";
    tmp(46644) := x"08e0";
    tmp(46645) := x"08e0";
    tmp(46646) := x"08e0";
    tmp(46647) := x"08e0";
    tmp(46648) := x"08e0";
    tmp(46649) := x"0900";
    tmp(46650) := x"0900";
    tmp(46651) := x"0900";
    tmp(46652) := x"0900";
    tmp(46653) := x"0900";
    tmp(46654) := x"0900";
    tmp(46655) := x"0900";
    tmp(46656) := x"0900";
    tmp(46657) := x"0920";
    tmp(46658) := x"0920";
    tmp(46659) := x"08a0";
    tmp(46660) := x"0020";
    tmp(46661) := x"0020";
    tmp(46662) := x"0021";
    tmp(46663) := x"0861";
    tmp(46664) := x"1082";
    tmp(46665) := x"0861";
    tmp(46666) := x"1082";
    tmp(46667) := x"0841";
    tmp(46668) := x"0841";
    tmp(46669) := x"0861";
    tmp(46670) := x"1082";
    tmp(46671) := x"1081";
    tmp(46672) := x"18c2";
    tmp(46673) := x"20e3";
    tmp(46674) := x"18c2";
    tmp(46675) := x"1061";
    tmp(46676) := x"0841";
    tmp(46677) := x"0841";
    tmp(46678) := x"0821";
    tmp(46679) := x"0861";
    tmp(46680) := x"0862";
    tmp(46681) := x"0841";
    tmp(46682) := x"0861";
    tmp(46683) := x"0861";
    tmp(46684) := x"0841";
    tmp(46685) := x"0861";
    tmp(46686) := x"0841";
    tmp(46687) := x"0841";
    tmp(46688) := x"0841";
    tmp(46689) := x"0841";
    tmp(46690) := x"0821";
    tmp(46691) := x"0820";
    tmp(46692) := x"0820";
    tmp(46693) := x"0821";
    tmp(46694) := x"0821";
    tmp(46695) := x"0821";
    tmp(46696) := x"0020";
    tmp(46697) := x"0000";
    tmp(46698) := x"0000";
    tmp(46699) := x"0000";
    tmp(46700) := x"0000";
    tmp(46701) := x"0000";
    tmp(46702) := x"0000";
    tmp(46703) := x"0020";
    tmp(46704) := x"0020";
    tmp(46705) := x"0821";
    tmp(46706) := x"0020";
    tmp(46707) := x"0000";
    tmp(46708) := x"0000";
    tmp(46709) := x"2081";
    tmp(46710) := x"3041";
    tmp(46711) := x"1800";
    tmp(46712) := x"1800";
    tmp(46713) := x"1800";
    tmp(46714) := x"1800";
    tmp(46715) := x"1800";
    tmp(46716) := x"2800";
    tmp(46717) := x"4861";
    tmp(46718) := x"3020";
    tmp(46719) := x"2820";
    tmp(46720) := x"68c3";
    tmp(46721) := x"50a2";
    tmp(46722) := x"2000";
    tmp(46723) := x"1800";
    tmp(46724) := x"2000";
    tmp(46725) := x"2000";
    tmp(46726) := x"3000";
    tmp(46727) := x"3800";
    tmp(46728) := x"3800";
    tmp(46729) := x"4800";
    tmp(46730) := x"5000";
    tmp(46731) := x"6000";
    tmp(46732) := x"7000";
    tmp(46733) := x"8800";
    tmp(46734) := x"8800";
    tmp(46735) := x"8800";
    tmp(46736) := x"9820";
    tmp(46737) := x"b020";
    tmp(46738) := x"a820";
    tmp(46739) := x"c020";
    tmp(46740) := x"c020";
    tmp(46741) := x"c020";
    tmp(46742) := x"d020";
    tmp(46743) := x"d820";
    tmp(46744) := x"f861";
    tmp(46745) := x"c861";
    tmp(46746) := x"4061";
    tmp(46747) := x"1040";
    tmp(46748) := x"1040";
    tmp(46749) := x"1040";
    tmp(46750) := x"0840";
    tmp(46751) := x"0840";
    tmp(46752) := x"0840";
    tmp(46753) := x"0840";
    tmp(46754) := x"0840";
    tmp(46755) := x"0840";
    tmp(46756) := x"0840";
    tmp(46757) := x"001f";
    tmp(46758) := x"001f";
    tmp(46759) := x"001f";
    tmp(46760) := x"001f";
    tmp(46761) := x"001f";
    tmp(46762) := x"001f";
    tmp(46763) := x"001f";
    tmp(46764) := x"001f";
    tmp(46765) := x"001f";
    tmp(46766) := x"001f";
    tmp(46767) := x"001f";
    tmp(46768) := x"001f";
    tmp(46769) := x"001f";
    tmp(46770) := x"001f";
    tmp(46771) := x"001f";
    tmp(46772) := x"001f";
    tmp(46773) := x"001f";
    tmp(46774) := x"001f";
    tmp(46775) := x"001f";
    tmp(46776) := x"001f";
    tmp(46777) := x"001f";
    tmp(46778) := x"001f";
    tmp(46779) := x"001f";
    tmp(46780) := x"001f";
    tmp(46781) := x"001f";
    tmp(46782) := x"001f";
    tmp(46783) := x"001f";
    tmp(46784) := x"001f";
    tmp(46785) := x"001f";
    tmp(46786) := x"001f";
    tmp(46787) := x"001f";
    tmp(46788) := x"001f";
    tmp(46789) := x"001f";
    tmp(46790) := x"001f";
    tmp(46791) := x"001f";
    tmp(46792) := x"001f";
    tmp(46793) := x"001f";
    tmp(46794) := x"001f";
    tmp(46795) := x"001f";
    tmp(46796) := x"001f";
    tmp(46797) := x"1040";
    tmp(46798) := x"0840";
    tmp(46799) := x"0840";
    tmp(46800) := x"0020";
    tmp(46801) := x"08c0";
    tmp(46802) := x"08c1";
    tmp(46803) := x"08c1";
    tmp(46804) := x"08c1";
    tmp(46805) := x"08c1";
    tmp(46806) := x"08e1";
    tmp(46807) := x"10e1";
    tmp(46808) := x"1101";
    tmp(46809) := x"1101";
    tmp(46810) := x"1101";
    tmp(46811) := x"10e1";
    tmp(46812) := x"10e1";
    tmp(46813) := x"10e1";
    tmp(46814) := x"10e1";
    tmp(46815) := x"10e1";
    tmp(46816) := x"10c1";
    tmp(46817) := x"10e1";
    tmp(46818) := x"10c1";
    tmp(46819) := x"10c1";
    tmp(46820) := x"10c1";
    tmp(46821) := x"10a1";
    tmp(46822) := x"10a1";
    tmp(46823) := x"08a1";
    tmp(46824) := x"08a1";
    tmp(46825) := x"08a1";
    tmp(46826) := x"08a1";
    tmp(46827) := x"10a1";
    tmp(46828) := x"10a1";
    tmp(46829) := x"10a1";
    tmp(46830) := x"10a1";
    tmp(46831) := x"10a1";
    tmp(46832) := x"10a1";
    tmp(46833) := x"1081";
    tmp(46834) := x"1081";
    tmp(46835) := x"1081";
    tmp(46836) := x"1081";
    tmp(46837) := x"0881";
    tmp(46838) := x"0861";
    tmp(46839) := x"0861";
    tmp(46840) := x"0861";
    tmp(46841) := x"0861";
    tmp(46842) := x"0861";
    tmp(46843) := x"0860";
    tmp(46844) := x"0860";
    tmp(46845) := x"0860";
    tmp(46846) := x"0860";
    tmp(46847) := x"0860";
    tmp(46848) := x"0860";
    tmp(46849) := x"0880";
    tmp(46850) := x"0880";
    tmp(46851) := x"0880";
    tmp(46852) := x"08a0";
    tmp(46853) := x"08a0";
    tmp(46854) := x"08a0";
    tmp(46855) := x"08a0";
    tmp(46856) := x"08a0";
    tmp(46857) := x"08c0";
    tmp(46858) := x"08c0";
    tmp(46859) := x"08c0";
    tmp(46860) := x"08c0";
    tmp(46861) := x"08c0";
    tmp(46862) := x"08c0";
    tmp(46863) := x"08c0";
    tmp(46864) := x"08e0";
    tmp(46865) := x"08e0";
    tmp(46866) := x"08e0";
    tmp(46867) := x"08e0";
    tmp(46868) := x"08e0";
    tmp(46869) := x"08e0";
    tmp(46870) := x"08c0";
    tmp(46871) := x"08c0";
    tmp(46872) := x"08c0";
    tmp(46873) := x"08c0";
    tmp(46874) := x"08c0";
    tmp(46875) := x"08c0";
    tmp(46876) := x"08c0";
    tmp(46877) := x"08c0";
    tmp(46878) := x"08c0";
    tmp(46879) := x"08c0";
    tmp(46880) := x"08c0";
    tmp(46881) := x"08c0";
    tmp(46882) := x"08e0";
    tmp(46883) := x"08e0";
    tmp(46884) := x"08e0";
    tmp(46885) := x"08e0";
    tmp(46886) := x"08e0";
    tmp(46887) := x"08e0";
    tmp(46888) := x"08e0";
    tmp(46889) := x"08e0";
    tmp(46890) := x"08e0";
    tmp(46891) := x"0900";
    tmp(46892) := x"08e0";
    tmp(46893) := x"0900";
    tmp(46894) := x"0900";
    tmp(46895) := x"0900";
    tmp(46896) := x"0900";
    tmp(46897) := x"0920";
    tmp(46898) := x"0900";
    tmp(46899) := x"0040";
    tmp(46900) := x"0000";
    tmp(46901) := x"0020";
    tmp(46902) := x"0021";
    tmp(46903) := x"0841";
    tmp(46904) := x"0841";
    tmp(46905) := x"0841";
    tmp(46906) := x"0841";
    tmp(46907) := x"0820";
    tmp(46908) := x"0820";
    tmp(46909) := x"0861";
    tmp(46910) := x"0861";
    tmp(46911) := x"1060";
    tmp(46912) := x"1060";
    tmp(46913) := x"0840";
    tmp(46914) := x"0841";
    tmp(46915) := x"0820";
    tmp(46916) := x"0820";
    tmp(46917) := x"0841";
    tmp(46918) := x"0861";
    tmp(46919) := x"0841";
    tmp(46920) := x"0020";
    tmp(46921) := x"0020";
    tmp(46922) := x"0020";
    tmp(46923) := x"0020";
    tmp(46924) := x"0000";
    tmp(46925) := x"0000";
    tmp(46926) := x"0000";
    tmp(46927) := x"0000";
    tmp(46928) := x"0020";
    tmp(46929) := x"0000";
    tmp(46930) := x"0000";
    tmp(46931) := x"0000";
    tmp(46932) := x"0000";
    tmp(46933) := x"0000";
    tmp(46934) := x"0000";
    tmp(46935) := x"0000";
    tmp(46936) := x"0000";
    tmp(46937) := x"0000";
    tmp(46938) := x"0000";
    tmp(46939) := x"0000";
    tmp(46940) := x"0000";
    tmp(46941) := x"0000";
    tmp(46942) := x"0000";
    tmp(46943) := x"0000";
    tmp(46944) := x"0000";
    tmp(46945) := x"0000";
    tmp(46946) := x"0000";
    tmp(46947) := x"0000";
    tmp(46948) := x"0000";
    tmp(46949) := x"3881";
    tmp(46950) := x"1800";
    tmp(46951) := x"1800";
    tmp(46952) := x"2000";
    tmp(46953) := x"2000";
    tmp(46954) := x"2000";
    tmp(46955) := x"2000";
    tmp(46956) := x"4061";
    tmp(46957) := x"58a2";
    tmp(46958) := x"3841";
    tmp(46959) := x"5082";
    tmp(46960) := x"68e4";
    tmp(46961) := x"3841";
    tmp(46962) := x"1800";
    tmp(46963) := x"1000";
    tmp(46964) := x"1800";
    tmp(46965) := x"2000";
    tmp(46966) := x"2800";
    tmp(46967) := x"3000";
    tmp(46968) := x"4000";
    tmp(46969) := x"4000";
    tmp(46970) := x"5000";
    tmp(46971) := x"6000";
    tmp(46972) := x"7000";
    tmp(46973) := x"7800";
    tmp(46974) := x"8800";
    tmp(46975) := x"9020";
    tmp(46976) := x"9820";
    tmp(46977) := x"b020";
    tmp(46978) := x"a800";
    tmp(46979) := x"b820";
    tmp(46980) := x"c820";
    tmp(46981) := x"c820";
    tmp(46982) := x"d020";
    tmp(46983) := x"d020";
    tmp(46984) := x"e841";
    tmp(46985) := x"f061";
    tmp(46986) := x"8061";
    tmp(46987) := x"1840";
    tmp(46988) := x"1040";
    tmp(46989) := x"1040";
    tmp(46990) := x"0840";
    tmp(46991) := x"0840";
    tmp(46992) := x"0840";
    tmp(46993) := x"0840";
    tmp(46994) := x"0840";
    tmp(46995) := x"0840";
    tmp(46996) := x"0840";
    tmp(46997) := x"001f";
    tmp(46998) := x"001f";
    tmp(46999) := x"001f";
    tmp(47000) := x"001f";
    tmp(47001) := x"001f";
    tmp(47002) := x"001f";
    tmp(47003) := x"001f";
    tmp(47004) := x"001f";
    tmp(47005) := x"001f";
    tmp(47006) := x"001f";
    tmp(47007) := x"001f";
    tmp(47008) := x"001f";
    tmp(47009) := x"001f";
    tmp(47010) := x"001f";
    tmp(47011) := x"001f";
    tmp(47012) := x"001f";
    tmp(47013) := x"001f";
    tmp(47014) := x"001f";
    tmp(47015) := x"001f";
    tmp(47016) := x"001f";
    tmp(47017) := x"001f";
    tmp(47018) := x"001f";
    tmp(47019) := x"001f";
    tmp(47020) := x"001f";
    tmp(47021) := x"001f";
    tmp(47022) := x"001f";
    tmp(47023) := x"001f";
    tmp(47024) := x"001f";
    tmp(47025) := x"001f";
    tmp(47026) := x"001f";
    tmp(47027) := x"001f";
    tmp(47028) := x"001f";
    tmp(47029) := x"001f";
    tmp(47030) := x"001f";
    tmp(47031) := x"001f";
    tmp(47032) := x"001f";
    tmp(47033) := x"001f";
    tmp(47034) := x"001f";
    tmp(47035) := x"001f";
    tmp(47036) := x"001f";
    tmp(47037) := x"0840";
    tmp(47038) := x"0840";
    tmp(47039) := x"0840";
    tmp(47040) := x"0020";
    tmp(47041) := x"08e1";
    tmp(47042) := x"08c0";
    tmp(47043) := x"08c1";
    tmp(47044) := x"08e1";
    tmp(47045) := x"08e1";
    tmp(47046) := x"08e1";
    tmp(47047) := x"10e1";
    tmp(47048) := x"10e1";
    tmp(47049) := x"10e1";
    tmp(47050) := x"1101";
    tmp(47051) := x"1101";
    tmp(47052) := x"1101";
    tmp(47053) := x"1101";
    tmp(47054) := x"10e1";
    tmp(47055) := x"10e1";
    tmp(47056) := x"10e1";
    tmp(47057) := x"10e1";
    tmp(47058) := x"10e1";
    tmp(47059) := x"10e1";
    tmp(47060) := x"10c1";
    tmp(47061) := x"10c1";
    tmp(47062) := x"10c1";
    tmp(47063) := x"10a1";
    tmp(47064) := x"08a1";
    tmp(47065) := x"08a1";
    tmp(47066) := x"08a1";
    tmp(47067) := x"10a1";
    tmp(47068) := x"10a1";
    tmp(47069) := x"10a1";
    tmp(47070) := x"10a1";
    tmp(47071) := x"10a1";
    tmp(47072) := x"10a1";
    tmp(47073) := x"10a1";
    tmp(47074) := x"1081";
    tmp(47075) := x"1081";
    tmp(47076) := x"1081";
    tmp(47077) := x"1081";
    tmp(47078) := x"0861";
    tmp(47079) := x"0861";
    tmp(47080) := x"0861";
    tmp(47081) := x"0861";
    tmp(47082) := x"0861";
    tmp(47083) := x"0860";
    tmp(47084) := x"0861";
    tmp(47085) := x"0860";
    tmp(47086) := x"0860";
    tmp(47087) := x"0860";
    tmp(47088) := x"0860";
    tmp(47089) := x"0860";
    tmp(47090) := x"0860";
    tmp(47091) := x"0880";
    tmp(47092) := x"0880";
    tmp(47093) := x"08a0";
    tmp(47094) := x"08a0";
    tmp(47095) := x"08a0";
    tmp(47096) := x"08a0";
    tmp(47097) := x"08a0";
    tmp(47098) := x"08c0";
    tmp(47099) := x"08c0";
    tmp(47100) := x"08c0";
    tmp(47101) := x"08c0";
    tmp(47102) := x"08c0";
    tmp(47103) := x"08c0";
    tmp(47104) := x"08c0";
    tmp(47105) := x"08c0";
    tmp(47106) := x"08c0";
    tmp(47107) := x"08c0";
    tmp(47108) := x"08c0";
    tmp(47109) := x"08c0";
    tmp(47110) := x"08c0";
    tmp(47111) := x"08c0";
    tmp(47112) := x"08c0";
    tmp(47113) := x"08c0";
    tmp(47114) := x"08c0";
    tmp(47115) := x"08c0";
    tmp(47116) := x"08c0";
    tmp(47117) := x"08c0";
    tmp(47118) := x"08c0";
    tmp(47119) := x"08c0";
    tmp(47120) := x"08c0";
    tmp(47121) := x"08c0";
    tmp(47122) := x"08c0";
    tmp(47123) := x"08c0";
    tmp(47124) := x"08c0";
    tmp(47125) := x"08c0";
    tmp(47126) := x"08e0";
    tmp(47127) := x"08e0";
    tmp(47128) := x"08e0";
    tmp(47129) := x"08e0";
    tmp(47130) := x"08e0";
    tmp(47131) := x"08e0";
    tmp(47132) := x"08e0";
    tmp(47133) := x"08e0";
    tmp(47134) := x"08e0";
    tmp(47135) := x"0900";
    tmp(47136) := x"0900";
    tmp(47137) := x"0900";
    tmp(47138) := x"08a0";
    tmp(47139) := x"0020";
    tmp(47140) := x"0000";
    tmp(47141) := x"0000";
    tmp(47142) := x"0020";
    tmp(47143) := x"0020";
    tmp(47144) := x"0020";
    tmp(47145) := x"0020";
    tmp(47146) := x"0020";
    tmp(47147) := x"0840";
    tmp(47148) := x"0860";
    tmp(47149) := x"0880";
    tmp(47150) := x"0880";
    tmp(47151) := x"10a0";
    tmp(47152) := x"0840";
    tmp(47153) := x"0000";
    tmp(47154) := x"0841";
    tmp(47155) := x"0841";
    tmp(47156) := x"0020";
    tmp(47157) := x"0020";
    tmp(47158) := x"0820";
    tmp(47159) := x"0820";
    tmp(47160) := x"0020";
    tmp(47161) := x"0000";
    tmp(47162) := x"0000";
    tmp(47163) := x"0000";
    tmp(47164) := x"0000";
    tmp(47165) := x"0000";
    tmp(47166) := x"0000";
    tmp(47167) := x"0000";
    tmp(47168) := x"0000";
    tmp(47169) := x"0000";
    tmp(47170) := x"0000";
    tmp(47171) := x"0000";
    tmp(47172) := x"0000";
    tmp(47173) := x"0000";
    tmp(47174) := x"0000";
    tmp(47175) := x"0000";
    tmp(47176) := x"0000";
    tmp(47177) := x"0000";
    tmp(47178) := x"0000";
    tmp(47179) := x"0000";
    tmp(47180) := x"0000";
    tmp(47181) := x"0000";
    tmp(47182) := x"0000";
    tmp(47183) := x"0000";
    tmp(47184) := x"0000";
    tmp(47185) := x"0000";
    tmp(47186) := x"0000";
    tmp(47187) := x"0000";
    tmp(47188) := x"1841";
    tmp(47189) := x"2820";
    tmp(47190) := x"1800";
    tmp(47191) := x"2000";
    tmp(47192) := x"2800";
    tmp(47193) := x"3020";
    tmp(47194) := x"3020";
    tmp(47195) := x"2820";
    tmp(47196) := x"3841";
    tmp(47197) := x"5082";
    tmp(47198) := x"4862";
    tmp(47199) := x"68e4";
    tmp(47200) := x"8125";
    tmp(47201) := x"a986";
    tmp(47202) := x"68a3";
    tmp(47203) := x"3841";
    tmp(47204) := x"1800";
    tmp(47205) := x"1800";
    tmp(47206) := x"2800";
    tmp(47207) := x"3000";
    tmp(47208) := x"4000";
    tmp(47209) := x"4800";
    tmp(47210) := x"5000";
    tmp(47211) := x"6000";
    tmp(47212) := x"6800";
    tmp(47213) := x"7800";
    tmp(47214) := x"8800";
    tmp(47215) := x"9820";
    tmp(47216) := x"a020";
    tmp(47217) := x"a820";
    tmp(47218) := x"9800";
    tmp(47219) := x"b020";
    tmp(47220) := x"c020";
    tmp(47221) := x"c820";
    tmp(47222) := x"c820";
    tmp(47223) := x"d820";
    tmp(47224) := x"d820";
    tmp(47225) := x"f041";
    tmp(47226) := x"c061";
    tmp(47227) := x"3861";
    tmp(47228) := x"1040";
    tmp(47229) := x"1040";
    tmp(47230) := x"1040";
    tmp(47231) := x"0840";
    tmp(47232) := x"0840";
    tmp(47233) := x"0840";
    tmp(47234) := x"0840";
    tmp(47235) := x"0840";
    tmp(47236) := x"0840";
    tmp(47237) := x"001f";
    tmp(47238) := x"001f";
    tmp(47239) := x"001f";
    tmp(47240) := x"001f";
    tmp(47241) := x"001f";
    tmp(47242) := x"001f";
    tmp(47243) := x"001f";
    tmp(47244) := x"001f";
    tmp(47245) := x"001f";
    tmp(47246) := x"001f";
    tmp(47247) := x"001f";
    tmp(47248) := x"001f";
    tmp(47249) := x"001f";
    tmp(47250) := x"001f";
    tmp(47251) := x"001f";
    tmp(47252) := x"001f";
    tmp(47253) := x"001f";
    tmp(47254) := x"001f";
    tmp(47255) := x"001f";
    tmp(47256) := x"001f";
    tmp(47257) := x"001f";
    tmp(47258) := x"001f";
    tmp(47259) := x"001f";
    tmp(47260) := x"001f";
    tmp(47261) := x"001f";
    tmp(47262) := x"001f";
    tmp(47263) := x"001f";
    tmp(47264) := x"001f";
    tmp(47265) := x"001f";
    tmp(47266) := x"001f";
    tmp(47267) := x"001f";
    tmp(47268) := x"001f";
    tmp(47269) := x"001f";
    tmp(47270) := x"001f";
    tmp(47271) := x"001f";
    tmp(47272) := x"001f";
    tmp(47273) := x"001f";
    tmp(47274) := x"001f";
    tmp(47275) := x"001f";
    tmp(47276) := x"001f";
    tmp(47277) := x"0840";
    tmp(47278) := x"0840";
    tmp(47279) := x"0840";
    tmp(47280) := x"0020";
    tmp(47281) := x"08c0";
    tmp(47282) := x"08c0";
    tmp(47283) := x"08c1";
    tmp(47284) := x"08c1";
    tmp(47285) := x"08c1";
    tmp(47286) := x"08e1";
    tmp(47287) := x"08e1";
    tmp(47288) := x"10e1";
    tmp(47289) := x"1101";
    tmp(47290) := x"1101";
    tmp(47291) := x"1101";
    tmp(47292) := x"1101";
    tmp(47293) := x"1101";
    tmp(47294) := x"1101";
    tmp(47295) := x"10e1";
    tmp(47296) := x"10e1";
    tmp(47297) := x"10e1";
    tmp(47298) := x"10e1";
    tmp(47299) := x"10e1";
    tmp(47300) := x"10e1";
    tmp(47301) := x"10e1";
    tmp(47302) := x"10e1";
    tmp(47303) := x"10c1";
    tmp(47304) := x"10c1";
    tmp(47305) := x"10a1";
    tmp(47306) := x"10a1";
    tmp(47307) := x"10a1";
    tmp(47308) := x"10a1";
    tmp(47309) := x"10a1";
    tmp(47310) := x"10a1";
    tmp(47311) := x"10a1";
    tmp(47312) := x"10a1";
    tmp(47313) := x"10a1";
    tmp(47314) := x"10a1";
    tmp(47315) := x"1081";
    tmp(47316) := x"0881";
    tmp(47317) := x"0881";
    tmp(47318) := x"0861";
    tmp(47319) := x"0861";
    tmp(47320) := x"0861";
    tmp(47321) := x"0861";
    tmp(47322) := x"0861";
    tmp(47323) := x"0861";
    tmp(47324) := x"0861";
    tmp(47325) := x"0861";
    tmp(47326) := x"0861";
    tmp(47327) := x"0860";
    tmp(47328) := x"0860";
    tmp(47329) := x"0860";
    tmp(47330) := x"0860";
    tmp(47331) := x"0880";
    tmp(47332) := x"0880";
    tmp(47333) := x"0880";
    tmp(47334) := x"08a0";
    tmp(47335) := x"08a0";
    tmp(47336) := x"08a0";
    tmp(47337) := x"08a0";
    tmp(47338) := x"08a0";
    tmp(47339) := x"08a0";
    tmp(47340) := x"08c0";
    tmp(47341) := x"08c0";
    tmp(47342) := x"08c0";
    tmp(47343) := x"08c0";
    tmp(47344) := x"08c0";
    tmp(47345) := x"08c0";
    tmp(47346) := x"08c0";
    tmp(47347) := x"08c0";
    tmp(47348) := x"08c0";
    tmp(47349) := x"08c0";
    tmp(47350) := x"08c0";
    tmp(47351) := x"08c0";
    tmp(47352) := x"08a0";
    tmp(47353) := x"08c0";
    tmp(47354) := x"08c0";
    tmp(47355) := x"08c0";
    tmp(47356) := x"08c0";
    tmp(47357) := x"08c0";
    tmp(47358) := x"08c0";
    tmp(47359) := x"08c0";
    tmp(47360) := x"08c0";
    tmp(47361) := x"08c0";
    tmp(47362) := x"08c0";
    tmp(47363) := x"08c0";
    tmp(47364) := x"08c0";
    tmp(47365) := x"08c0";
    tmp(47366) := x"08c0";
    tmp(47367) := x"08c0";
    tmp(47368) := x"08c0";
    tmp(47369) := x"08e0";
    tmp(47370) := x"08c0";
    tmp(47371) := x"08e0";
    tmp(47372) := x"08e0";
    tmp(47373) := x"08e0";
    tmp(47374) := x"08e0";
    tmp(47375) := x"0900";
    tmp(47376) := x"0900";
    tmp(47377) := x"0900";
    tmp(47378) := x"0040";
    tmp(47379) := x"0000";
    tmp(47380) := x"0000";
    tmp(47381) := x"0000";
    tmp(47382) := x"0020";
    tmp(47383) := x"0000";
    tmp(47384) := x"0020";
    tmp(47385) := x"0840";
    tmp(47386) := x"0860";
    tmp(47387) := x"08a0";
    tmp(47388) := x"10a0";
    tmp(47389) := x"08a0";
    tmp(47390) := x"10a0";
    tmp(47391) := x"0860";
    tmp(47392) := x"0820";
    tmp(47393) := x"0000";
    tmp(47394) := x"0020";
    tmp(47395) := x"0841";
    tmp(47396) := x"0020";
    tmp(47397) := x"0000";
    tmp(47398) := x"0000";
    tmp(47399) := x"0020";
    tmp(47400) := x"0020";
    tmp(47401) := x"0000";
    tmp(47402) := x"0000";
    tmp(47403) := x"0000";
    tmp(47404) := x"0000";
    tmp(47405) := x"0000";
    tmp(47406) := x"0000";
    tmp(47407) := x"0000";
    tmp(47408) := x"0000";
    tmp(47409) := x"0000";
    tmp(47410) := x"0000";
    tmp(47411) := x"0000";
    tmp(47412) := x"0000";
    tmp(47413) := x"0000";
    tmp(47414) := x"0000";
    tmp(47415) := x"0000";
    tmp(47416) := x"0000";
    tmp(47417) := x"0000";
    tmp(47418) := x"0000";
    tmp(47419) := x"0000";
    tmp(47420) := x"0000";
    tmp(47421) := x"0000";
    tmp(47422) := x"0000";
    tmp(47423) := x"0000";
    tmp(47424) := x"0000";
    tmp(47425) := x"0000";
    tmp(47426) := x"0000";
    tmp(47427) := x"0820";
    tmp(47428) := x"3061";
    tmp(47429) := x"2000";
    tmp(47430) := x"2000";
    tmp(47431) := x"2800";
    tmp(47432) := x"4041";
    tmp(47433) := x"68e4";
    tmp(47434) := x"4861";
    tmp(47435) := x"2820";
    tmp(47436) := x"3021";
    tmp(47437) := x"5082";
    tmp(47438) := x"58a3";
    tmp(47439) := x"7925";
    tmp(47440) := x"70e4";
    tmp(47441) := x"5082";
    tmp(47442) := x"ca09";
    tmp(47443) := x"8925";
    tmp(47444) := x"2820";
    tmp(47445) := x"1800";
    tmp(47446) := x"2000";
    tmp(47447) := x"3000";
    tmp(47448) := x"4000";
    tmp(47449) := x"4800";
    tmp(47450) := x"5000";
    tmp(47451) := x"6000";
    tmp(47452) := x"6800";
    tmp(47453) := x"8000";
    tmp(47454) := x"8800";
    tmp(47455) := x"8800";
    tmp(47456) := x"a820";
    tmp(47457) := x"a020";
    tmp(47458) := x"9820";
    tmp(47459) := x"a820";
    tmp(47460) := x"b020";
    tmp(47461) := x"d020";
    tmp(47462) := x"d820";
    tmp(47463) := x"d820";
    tmp(47464) := x"d820";
    tmp(47465) := x"f041";
    tmp(47466) := x"d861";
    tmp(47467) := x"6861";
    tmp(47468) := x"1840";
    tmp(47469) := x"1040";
    tmp(47470) := x"1040";
    tmp(47471) := x"1040";
    tmp(47472) := x"1040";
    tmp(47473) := x"0840";
    tmp(47474) := x"0840";
    tmp(47475) := x"0840";
    tmp(47476) := x"0840";
    tmp(47477) := x"001f";
    tmp(47478) := x"001f";
    tmp(47479) := x"001f";
    tmp(47480) := x"001f";
    tmp(47481) := x"001f";
    tmp(47482) := x"001f";
    tmp(47483) := x"001f";
    tmp(47484) := x"001f";
    tmp(47485) := x"001f";
    tmp(47486) := x"001f";
    tmp(47487) := x"001f";
    tmp(47488) := x"001f";
    tmp(47489) := x"001f";
    tmp(47490) := x"001f";
    tmp(47491) := x"001f";
    tmp(47492) := x"001f";
    tmp(47493) := x"001f";
    tmp(47494) := x"001f";
    tmp(47495) := x"001f";
    tmp(47496) := x"001f";
    tmp(47497) := x"001f";
    tmp(47498) := x"001f";
    tmp(47499) := x"001f";
    tmp(47500) := x"001f";
    tmp(47501) := x"001f";
    tmp(47502) := x"001f";
    tmp(47503) := x"001f";
    tmp(47504) := x"001f";
    tmp(47505) := x"001f";
    tmp(47506) := x"001f";
    tmp(47507) := x"001f";
    tmp(47508) := x"001f";
    tmp(47509) := x"001f";
    tmp(47510) := x"001f";
    tmp(47511) := x"001f";
    tmp(47512) := x"001f";
    tmp(47513) := x"001f";
    tmp(47514) := x"001f";
    tmp(47515) := x"001f";
    tmp(47516) := x"001f";
    tmp(47517) := x"0840";
    tmp(47518) := x"0840";
    tmp(47519) := x"0840";
    tmp(47520) := x"0020";
    tmp(47521) := x"08c0";
    tmp(47522) := x"08c0";
    tmp(47523) := x"08c1";
    tmp(47524) := x"08c1";
    tmp(47525) := x"08e1";
    tmp(47526) := x"08e1";
    tmp(47527) := x"08e1";
    tmp(47528) := x"08e1";
    tmp(47529) := x"1101";
    tmp(47530) := x"1101";
    tmp(47531) := x"1101";
    tmp(47532) := x"1101";
    tmp(47533) := x"1101";
    tmp(47534) := x"1101";
    tmp(47535) := x"1101";
    tmp(47536) := x"10e1";
    tmp(47537) := x"1101";
    tmp(47538) := x"1101";
    tmp(47539) := x"10e1";
    tmp(47540) := x"10e1";
    tmp(47541) := x"10e1";
    tmp(47542) := x"10e1";
    tmp(47543) := x"10e1";
    tmp(47544) := x"10e1";
    tmp(47545) := x"10c1";
    tmp(47546) := x"10c1";
    tmp(47547) := x"10c1";
    tmp(47548) := x"10a1";
    tmp(47549) := x"10c1";
    tmp(47550) := x"10a1";
    tmp(47551) := x"10a1";
    tmp(47552) := x"10a1";
    tmp(47553) := x"10a1";
    tmp(47554) := x"10a1";
    tmp(47555) := x"10a1";
    tmp(47556) := x"0881";
    tmp(47557) := x"0881";
    tmp(47558) := x"0881";
    tmp(47559) := x"0861";
    tmp(47560) := x"0861";
    tmp(47561) := x"0861";
    tmp(47562) := x"0861";
    tmp(47563) := x"0861";
    tmp(47564) := x"0861";
    tmp(47565) := x"0860";
    tmp(47566) := x"0861";
    tmp(47567) := x"0860";
    tmp(47568) := x"0861";
    tmp(47569) := x"0861";
    tmp(47570) := x"0860";
    tmp(47571) := x"0860";
    tmp(47572) := x"0880";
    tmp(47573) := x"0880";
    tmp(47574) := x"0880";
    tmp(47575) := x"0880";
    tmp(47576) := x"0880";
    tmp(47577) := x"08a0";
    tmp(47578) := x"08a0";
    tmp(47579) := x"08a1";
    tmp(47580) := x"08a0";
    tmp(47581) := x"08a0";
    tmp(47582) := x"08a0";
    tmp(47583) := x"08a0";
    tmp(47584) := x"08a0";
    tmp(47585) := x"08a0";
    tmp(47586) := x"08a0";
    tmp(47587) := x"08a0";
    tmp(47588) := x"08a0";
    tmp(47589) := x"08a0";
    tmp(47590) := x"08a0";
    tmp(47591) := x"08a0";
    tmp(47592) := x"08a0";
    tmp(47593) := x"08a0";
    tmp(47594) := x"08a0";
    tmp(47595) := x"08a0";
    tmp(47596) := x"08a0";
    tmp(47597) := x"08a0";
    tmp(47598) := x"08a0";
    tmp(47599) := x"08a0";
    tmp(47600) := x"08a0";
    tmp(47601) := x"08a0";
    tmp(47602) := x"08c0";
    tmp(47603) := x"08c0";
    tmp(47604) := x"08c0";
    tmp(47605) := x"08c0";
    tmp(47606) := x"08c0";
    tmp(47607) := x"08c0";
    tmp(47608) := x"08c0";
    tmp(47609) := x"08c0";
    tmp(47610) := x"08c0";
    tmp(47611) := x"08c0";
    tmp(47612) := x"08c0";
    tmp(47613) := x"08c0";
    tmp(47614) := x"08e0";
    tmp(47615) := x"08e0";
    tmp(47616) := x"08e0";
    tmp(47617) := x"08a0";
    tmp(47618) := x"0020";
    tmp(47619) := x"0000";
    tmp(47620) := x"0000";
    tmp(47621) := x"0000";
    tmp(47622) := x"0020";
    tmp(47623) := x"0840";
    tmp(47624) := x"0880";
    tmp(47625) := x"08a0";
    tmp(47626) := x"10c0";
    tmp(47627) := x"10a0";
    tmp(47628) := x"08a0";
    tmp(47629) := x"10a0";
    tmp(47630) := x"10a0";
    tmp(47631) := x"0860";
    tmp(47632) := x"0840";
    tmp(47633) := x"0000";
    tmp(47634) := x"0020";
    tmp(47635) := x"0841";
    tmp(47636) := x"0000";
    tmp(47637) := x"0000";
    tmp(47638) := x"0000";
    tmp(47639) := x"0000";
    tmp(47640) := x"0000";
    tmp(47641) := x"0000";
    tmp(47642) := x"0000";
    tmp(47643) := x"0000";
    tmp(47644) := x"0000";
    tmp(47645) := x"0000";
    tmp(47646) := x"0000";
    tmp(47647) := x"0000";
    tmp(47648) := x"0000";
    tmp(47649) := x"0000";
    tmp(47650) := x"0000";
    tmp(47651) := x"0000";
    tmp(47652) := x"0000";
    tmp(47653) := x"0000";
    tmp(47654) := x"0000";
    tmp(47655) := x"0000";
    tmp(47656) := x"0000";
    tmp(47657) := x"0000";
    tmp(47658) := x"0000";
    tmp(47659) := x"0000";
    tmp(47660) := x"0000";
    tmp(47661) := x"0000";
    tmp(47662) := x"0000";
    tmp(47663) := x"0000";
    tmp(47664) := x"0000";
    tmp(47665) := x"0000";
    tmp(47666) := x"0000";
    tmp(47667) := x"3081";
    tmp(47668) := x"2820";
    tmp(47669) := x"2000";
    tmp(47670) := x"4021";
    tmp(47671) := x"5862";
    tmp(47672) := x"70e4";
    tmp(47673) := x"7946";
    tmp(47674) := x"50a3";
    tmp(47675) := x"2820";
    tmp(47676) := x"2820";
    tmp(47677) := x"60a3";
    tmp(47678) := x"99a7";
    tmp(47679) := x"a9e9";
    tmp(47680) := x"68e4";
    tmp(47681) := x"5041";
    tmp(47682) := x"6082";
    tmp(47683) := x"68a2";
    tmp(47684) := x"2000";
    tmp(47685) := x"2000";
    tmp(47686) := x"2000";
    tmp(47687) := x"2800";
    tmp(47688) := x"3000";
    tmp(47689) := x"4000";
    tmp(47690) := x"4800";
    tmp(47691) := x"6000";
    tmp(47692) := x"7000";
    tmp(47693) := x"7800";
    tmp(47694) := x"8800";
    tmp(47695) := x"8800";
    tmp(47696) := x"9000";
    tmp(47697) := x"a020";
    tmp(47698) := x"b020";
    tmp(47699) := x"b020";
    tmp(47700) := x"c820";
    tmp(47701) := x"d820";
    tmp(47702) := x"c820";
    tmp(47703) := x"e020";
    tmp(47704) := x"e820";
    tmp(47705) := x"e840";
    tmp(47706) := x"d040";
    tmp(47707) := x"9061";
    tmp(47708) := x"2840";
    tmp(47709) := x"1040";
    tmp(47710) := x"1040";
    tmp(47711) := x"1040";
    tmp(47712) := x"1040";
    tmp(47713) := x"0840";
    tmp(47714) := x"0840";
    tmp(47715) := x"0840";
    tmp(47716) := x"0840";
    tmp(47717) := x"001f";
    tmp(47718) := x"001f";
    tmp(47719) := x"001f";
    tmp(47720) := x"001f";
    tmp(47721) := x"001f";
    tmp(47722) := x"001f";
    tmp(47723) := x"001f";
    tmp(47724) := x"001f";
    tmp(47725) := x"001f";
    tmp(47726) := x"001f";
    tmp(47727) := x"001f";
    tmp(47728) := x"001f";
    tmp(47729) := x"001f";
    tmp(47730) := x"001f";
    tmp(47731) := x"001f";
    tmp(47732) := x"001f";
    tmp(47733) := x"001f";
    tmp(47734) := x"001f";
    tmp(47735) := x"001f";
    tmp(47736) := x"001f";
    tmp(47737) := x"001f";
    tmp(47738) := x"001f";
    tmp(47739) := x"001f";
    tmp(47740) := x"001f";
    tmp(47741) := x"001f";
    tmp(47742) := x"001f";
    tmp(47743) := x"001f";
    tmp(47744) := x"001f";
    tmp(47745) := x"001f";
    tmp(47746) := x"001f";
    tmp(47747) := x"001f";
    tmp(47748) := x"001f";
    tmp(47749) := x"001f";
    tmp(47750) := x"001f";
    tmp(47751) := x"001f";
    tmp(47752) := x"001f";
    tmp(47753) := x"001f";
    tmp(47754) := x"001f";
    tmp(47755) := x"001f";
    tmp(47756) := x"001f";
    tmp(47757) := x"0840";
    tmp(47758) := x"0840";
    tmp(47759) := x"0840";
    tmp(47760) := x"0000";
    tmp(47761) := x"08c0";
    tmp(47762) := x"08c0";
    tmp(47763) := x"08c1";
    tmp(47764) := x"08c1";
    tmp(47765) := x"08c1";
    tmp(47766) := x"08e1";
    tmp(47767) := x"08e1";
    tmp(47768) := x"08e1";
    tmp(47769) := x"10e1";
    tmp(47770) := x"1101";
    tmp(47771) := x"1101";
    tmp(47772) := x"1101";
    tmp(47773) := x"1101";
    tmp(47774) := x"1101";
    tmp(47775) := x"10e1";
    tmp(47776) := x"1101";
    tmp(47777) := x"10e1";
    tmp(47778) := x"1101";
    tmp(47779) := x"1101";
    tmp(47780) := x"1101";
    tmp(47781) := x"1101";
    tmp(47782) := x"1101";
    tmp(47783) := x"10e1";
    tmp(47784) := x"1101";
    tmp(47785) := x"10e1";
    tmp(47786) := x"10e1";
    tmp(47787) := x"10e1";
    tmp(47788) := x"10c1";
    tmp(47789) := x"10c1";
    tmp(47790) := x"10c1";
    tmp(47791) := x"10c1";
    tmp(47792) := x"10a1";
    tmp(47793) := x"10a1";
    tmp(47794) := x"08a1";
    tmp(47795) := x"08a1";
    tmp(47796) := x"0881";
    tmp(47797) := x"0881";
    tmp(47798) := x"0881";
    tmp(47799) := x"0881";
    tmp(47800) := x"0861";
    tmp(47801) := x"0861";
    tmp(47802) := x"0861";
    tmp(47803) := x"0861";
    tmp(47804) := x"0861";
    tmp(47805) := x"0861";
    tmp(47806) := x"0861";
    tmp(47807) := x"0861";
    tmp(47808) := x"0861";
    tmp(47809) := x"0861";
    tmp(47810) := x"0861";
    tmp(47811) := x"0861";
    tmp(47812) := x"0860";
    tmp(47813) := x"0881";
    tmp(47814) := x"0881";
    tmp(47815) := x"0881";
    tmp(47816) := x"0881";
    tmp(47817) := x"08a1";
    tmp(47818) := x"08a0";
    tmp(47819) := x"08a1";
    tmp(47820) := x"08a0";
    tmp(47821) := x"08a0";
    tmp(47822) := x"08a0";
    tmp(47823) := x"08a0";
    tmp(47824) := x"08a0";
    tmp(47825) := x"08a0";
    tmp(47826) := x"08a0";
    tmp(47827) := x"08a0";
    tmp(47828) := x"08a0";
    tmp(47829) := x"08a0";
    tmp(47830) := x"08a0";
    tmp(47831) := x"08a0";
    tmp(47832) := x"08a0";
    tmp(47833) := x"08a0";
    tmp(47834) := x"08a0";
    tmp(47835) := x"08a0";
    tmp(47836) := x"08a0";
    tmp(47837) := x"08a0";
    tmp(47838) := x"08a0";
    tmp(47839) := x"08a0";
    tmp(47840) := x"08a0";
    tmp(47841) := x"08a0";
    tmp(47842) := x"08a0";
    tmp(47843) := x"08a0";
    tmp(47844) := x"08a0";
    tmp(47845) := x"08a0";
    tmp(47846) := x"08c0";
    tmp(47847) := x"08c0";
    tmp(47848) := x"08c0";
    tmp(47849) := x"08c0";
    tmp(47850) := x"08c0";
    tmp(47851) := x"08c0";
    tmp(47852) := x"08c0";
    tmp(47853) := x"08c0";
    tmp(47854) := x"08c0";
    tmp(47855) := x"08c0";
    tmp(47856) := x"08e0";
    tmp(47857) := x"0840";
    tmp(47858) := x"0000";
    tmp(47859) := x"0000";
    tmp(47860) := x"0000";
    tmp(47861) := x"0020";
    tmp(47862) := x"0880";
    tmp(47863) := x"10c0";
    tmp(47864) := x"10c0";
    tmp(47865) := x"08c0";
    tmp(47866) := x"10c0";
    tmp(47867) := x"10a0";
    tmp(47868) := x"08a0";
    tmp(47869) := x"10a0";
    tmp(47870) := x"1080";
    tmp(47871) := x"10a0";
    tmp(47872) := x"0860";
    tmp(47873) := x"0000";
    tmp(47874) := x"0820";
    tmp(47875) := x"1081";
    tmp(47876) := x"0000";
    tmp(47877) := x"0000";
    tmp(47878) := x"0000";
    tmp(47879) := x"0000";
    tmp(47880) := x"0000";
    tmp(47881) := x"0000";
    tmp(47882) := x"0000";
    tmp(47883) := x"0000";
    tmp(47884) := x"0000";
    tmp(47885) := x"0000";
    tmp(47886) := x"0000";
    tmp(47887) := x"0000";
    tmp(47888) := x"0000";
    tmp(47889) := x"0000";
    tmp(47890) := x"0000";
    tmp(47891) := x"0000";
    tmp(47892) := x"0000";
    tmp(47893) := x"0000";
    tmp(47894) := x"0000";
    tmp(47895) := x"0000";
    tmp(47896) := x"0000";
    tmp(47897) := x"0000";
    tmp(47898) := x"0000";
    tmp(47899) := x"0000";
    tmp(47900) := x"0000";
    tmp(47901) := x"0000";
    tmp(47902) := x"0000";
    tmp(47903) := x"0000";
    tmp(47904) := x"0000";
    tmp(47905) := x"0000";
    tmp(47906) := x"4104";
    tmp(47907) := x"4881";
    tmp(47908) := x"2800";
    tmp(47909) := x"3000";
    tmp(47910) := x"5882";
    tmp(47911) := x"60c3";
    tmp(47912) := x"60c4";
    tmp(47913) := x"99e9";
    tmp(47914) := x"8187";
    tmp(47915) := x"5082";
    tmp(47916) := x"5062";
    tmp(47917) := x"9146";
    tmp(47918) := x"8125";
    tmp(47919) := x"5082";
    tmp(47920) := x"78e4";
    tmp(47921) := x"c1c7";
    tmp(47922) := x"b9e8";
    tmp(47923) := x"c1c7";
    tmp(47924) := x"80c3";
    tmp(47925) := x"5041";
    tmp(47926) := x"2000";
    tmp(47927) := x"2000";
    tmp(47928) := x"2800";
    tmp(47929) := x"3800";
    tmp(47930) := x"4000";
    tmp(47931) := x"5800";
    tmp(47932) := x"7000";
    tmp(47933) := x"7800";
    tmp(47934) := x"8000";
    tmp(47935) := x"9020";
    tmp(47936) := x"8800";
    tmp(47937) := x"a020";
    tmp(47938) := x"b020";
    tmp(47939) := x"c020";
    tmp(47940) := x"c020";
    tmp(47941) := x"d020";
    tmp(47942) := x"e020";
    tmp(47943) := x"e020";
    tmp(47944) := x"f020";
    tmp(47945) := x"e020";
    tmp(47946) := x"d020";
    tmp(47947) := x"b861";
    tmp(47948) := x"3841";
    tmp(47949) := x"1040";
    tmp(47950) := x"1040";
    tmp(47951) := x"1040";
    tmp(47952) := x"0840";
    tmp(47953) := x"0840";
    tmp(47954) := x"0840";
    tmp(47955) := x"0840";
    tmp(47956) := x"0840";
    tmp(47957) := x"001f";
    tmp(47958) := x"001f";
    tmp(47959) := x"001f";
    tmp(47960) := x"001f";
    tmp(47961) := x"001f";
    tmp(47962) := x"001f";
    tmp(47963) := x"001f";
    tmp(47964) := x"001f";
    tmp(47965) := x"001f";
    tmp(47966) := x"001f";
    tmp(47967) := x"001f";
    tmp(47968) := x"001f";
    tmp(47969) := x"001f";
    tmp(47970) := x"001f";
    tmp(47971) := x"001f";
    tmp(47972) := x"001f";
    tmp(47973) := x"001f";
    tmp(47974) := x"001f";
    tmp(47975) := x"001f";
    tmp(47976) := x"001f";
    tmp(47977) := x"001f";
    tmp(47978) := x"001f";
    tmp(47979) := x"001f";
    tmp(47980) := x"001f";
    tmp(47981) := x"001f";
    tmp(47982) := x"001f";
    tmp(47983) := x"001f";
    tmp(47984) := x"001f";
    tmp(47985) := x"001f";
    tmp(47986) := x"001f";
    tmp(47987) := x"001f";
    tmp(47988) := x"001f";
    tmp(47989) := x"001f";
    tmp(47990) := x"001f";
    tmp(47991) := x"001f";
    tmp(47992) := x"001f";
    tmp(47993) := x"001f";
    tmp(47994) := x"001f";
    tmp(47995) := x"001f";
    tmp(47996) := x"001f";
    tmp(47997) := x"0840";
    tmp(47998) := x"0840";
    tmp(47999) := x"0840";
    tmp(48000) := x"0020";
    tmp(48001) := x"08c0";
    tmp(48002) := x"08c0";
    tmp(48003) := x"08e1";
    tmp(48004) := x"08e1";
    tmp(48005) := x"08e1";
    tmp(48006) := x"08e1";
    tmp(48007) := x"08e1";
    tmp(48008) := x"08e1";
    tmp(48009) := x"08e1";
    tmp(48010) := x"10e1";
    tmp(48011) := x"1101";
    tmp(48012) := x"1101";
    tmp(48013) := x"1101";
    tmp(48014) := x"1101";
    tmp(48015) := x"1101";
    tmp(48016) := x"1101";
    tmp(48017) := x"1101";
    tmp(48018) := x"1101";
    tmp(48019) := x"1101";
    tmp(48020) := x"1101";
    tmp(48021) := x"1101";
    tmp(48022) := x"1101";
    tmp(48023) := x"1101";
    tmp(48024) := x"1101";
    tmp(48025) := x"1101";
    tmp(48026) := x"1101";
    tmp(48027) := x"1101";
    tmp(48028) := x"10e1";
    tmp(48029) := x"10e1";
    tmp(48030) := x"10e1";
    tmp(48031) := x"10c1";
    tmp(48032) := x"10c1";
    tmp(48033) := x"10c1";
    tmp(48034) := x"08a1";
    tmp(48035) := x"08a1";
    tmp(48036) := x"0881";
    tmp(48037) := x"0881";
    tmp(48038) := x"0881";
    tmp(48039) := x"0881";
    tmp(48040) := x"0881";
    tmp(48041) := x"0861";
    tmp(48042) := x"0861";
    tmp(48043) := x"0861";
    tmp(48044) := x"0861";
    tmp(48045) := x"0861";
    tmp(48046) := x"0860";
    tmp(48047) := x"0861";
    tmp(48048) := x"0861";
    tmp(48049) := x"0860";
    tmp(48050) := x"0861";
    tmp(48051) := x"0861";
    tmp(48052) := x"0861";
    tmp(48053) := x"0861";
    tmp(48054) := x"0861";
    tmp(48055) := x"0881";
    tmp(48056) := x"0881";
    tmp(48057) := x"0881";
    tmp(48058) := x"0881";
    tmp(48059) := x"0881";
    tmp(48060) := x"08a1";
    tmp(48061) := x"08a1";
    tmp(48062) := x"08a1";
    tmp(48063) := x"08a1";
    tmp(48064) := x"08a1";
    tmp(48065) := x"08a1";
    tmp(48066) := x"08a1";
    tmp(48067) := x"08a1";
    tmp(48068) := x"08a1";
    tmp(48069) := x"08a1";
    tmp(48070) := x"08a1";
    tmp(48071) := x"08a1";
    tmp(48072) := x"08a1";
    tmp(48073) := x"08a0";
    tmp(48074) := x"08a0";
    tmp(48075) := x"08a0";
    tmp(48076) := x"08a0";
    tmp(48077) := x"08a0";
    tmp(48078) := x"08a0";
    tmp(48079) := x"08a0";
    tmp(48080) := x"08a0";
    tmp(48081) := x"08a0";
    tmp(48082) := x"08a0";
    tmp(48083) := x"08a0";
    tmp(48084) := x"08a0";
    tmp(48085) := x"08a0";
    tmp(48086) := x"08a0";
    tmp(48087) := x"08a0";
    tmp(48088) := x"08a0";
    tmp(48089) := x"08c0";
    tmp(48090) := x"08a0";
    tmp(48091) := x"08a0";
    tmp(48092) := x"08c0";
    tmp(48093) := x"08c0";
    tmp(48094) := x"08c0";
    tmp(48095) := x"08c0";
    tmp(48096) := x"08c0";
    tmp(48097) := x"0020";
    tmp(48098) := x"0000";
    tmp(48099) := x"0000";
    tmp(48100) := x"0020";
    tmp(48101) := x"08a0";
    tmp(48102) := x"10c0";
    tmp(48103) := x"10c0";
    tmp(48104) := x"10c0";
    tmp(48105) := x"10a0";
    tmp(48106) := x"10a0";
    tmp(48107) := x"10a0";
    tmp(48108) := x"10a0";
    tmp(48109) := x"0880";
    tmp(48110) := x"1080";
    tmp(48111) := x"1080";
    tmp(48112) := x"0840";
    tmp(48113) := x"0000";
    tmp(48114) := x"0000";
    tmp(48115) := x"0861";
    tmp(48116) := x"0020";
    tmp(48117) := x"0000";
    tmp(48118) := x"0000";
    tmp(48119) := x"0000";
    tmp(48120) := x"0000";
    tmp(48121) := x"0000";
    tmp(48122) := x"0000";
    tmp(48123) := x"0000";
    tmp(48124) := x"0000";
    tmp(48125) := x"0000";
    tmp(48126) := x"0000";
    tmp(48127) := x"0021";
    tmp(48128) := x"0020";
    tmp(48129) := x"0000";
    tmp(48130) := x"0000";
    tmp(48131) := x"0000";
    tmp(48132) := x"0000";
    tmp(48133) := x"0000";
    tmp(48134) := x"0000";
    tmp(48135) := x"0000";
    tmp(48136) := x"0000";
    tmp(48137) := x"0000";
    tmp(48138) := x"0000";
    tmp(48139) := x"0000";
    tmp(48140) := x"0000";
    tmp(48141) := x"0020";
    tmp(48142) := x"0000";
    tmp(48143) := x"0000";
    tmp(48144) := x"0000";
    tmp(48145) := x"4124";
    tmp(48146) := x"cb6d";
    tmp(48147) := x"70c3";
    tmp(48148) := x"3000";
    tmp(48149) := x"3020";
    tmp(48150) := x"3821";
    tmp(48151) := x"58a2";
    tmp(48152) := x"7104";
    tmp(48153) := x"89c8";
    tmp(48154) := x"99e9";
    tmp(48155) := x"7104";
    tmp(48156) := x"b208";
    tmp(48157) := x"e32e";
    tmp(48158) := x"e38f";
    tmp(48159) := x"8966";
    tmp(48160) := x"5882";
    tmp(48161) := x"4041";
    tmp(48162) := x"9125";
    tmp(48163) := x"ca08";
    tmp(48164) := x"da6a";
    tmp(48165) := x"5041";
    tmp(48166) := x"3820";
    tmp(48167) := x"2800";
    tmp(48168) := x"2800";
    tmp(48169) := x"3000";
    tmp(48170) := x"3800";
    tmp(48171) := x"5000";
    tmp(48172) := x"6800";
    tmp(48173) := x"7800";
    tmp(48174) := x"8000";
    tmp(48175) := x"8800";
    tmp(48176) := x"9820";
    tmp(48177) := x"a020";
    tmp(48178) := x"b020";
    tmp(48179) := x"c020";
    tmp(48180) := x"d820";
    tmp(48181) := x"c820";
    tmp(48182) := x"d020";
    tmp(48183) := x"d820";
    tmp(48184) := x"f040";
    tmp(48185) := x"e820";
    tmp(48186) := x"d020";
    tmp(48187) := x"c041";
    tmp(48188) := x"5061";
    tmp(48189) := x"1040";
    tmp(48190) := x"1040";
    tmp(48191) := x"0840";
    tmp(48192) := x"0840";
    tmp(48193) := x"0840";
    tmp(48194) := x"0840";
    tmp(48195) := x"0840";
    tmp(48196) := x"0840";
    tmp(48197) := x"001f";
    tmp(48198) := x"001f";
    tmp(48199) := x"001f";
    tmp(48200) := x"001f";
    tmp(48201) := x"001f";
    tmp(48202) := x"001f";
    tmp(48203) := x"001f";
    tmp(48204) := x"001f";
    tmp(48205) := x"001f";
    tmp(48206) := x"001f";
    tmp(48207) := x"001f";
    tmp(48208) := x"001f";
    tmp(48209) := x"001f";
    tmp(48210) := x"001f";
    tmp(48211) := x"001f";
    tmp(48212) := x"001f";
    tmp(48213) := x"001f";
    tmp(48214) := x"001f";
    tmp(48215) := x"001f";
    tmp(48216) := x"001f";
    tmp(48217) := x"001f";
    tmp(48218) := x"001f";
    tmp(48219) := x"001f";
    tmp(48220) := x"001f";
    tmp(48221) := x"001f";
    tmp(48222) := x"001f";
    tmp(48223) := x"001f";
    tmp(48224) := x"001f";
    tmp(48225) := x"001f";
    tmp(48226) := x"001f";
    tmp(48227) := x"001f";
    tmp(48228) := x"001f";
    tmp(48229) := x"001f";
    tmp(48230) := x"001f";
    tmp(48231) := x"001f";
    tmp(48232) := x"001f";
    tmp(48233) := x"001f";
    tmp(48234) := x"001f";
    tmp(48235) := x"001f";
    tmp(48236) := x"001f";
    tmp(48237) := x"0840";
    tmp(48238) := x"0840";
    tmp(48239) := x"0840";
    tmp(48240) := x"0020";
    tmp(48241) := x"08e1";
    tmp(48242) := x"08c1";
    tmp(48243) := x"08e1";
    tmp(48244) := x"08e1";
    tmp(48245) := x"08e1";
    tmp(48246) := x"08e1";
    tmp(48247) := x"08e1";
    tmp(48248) := x"08c1";
    tmp(48249) := x"08e1";
    tmp(48250) := x"08c1";
    tmp(48251) := x"10e1";
    tmp(48252) := x"10e1";
    tmp(48253) := x"1101";
    tmp(48254) := x"1101";
    tmp(48255) := x"1101";
    tmp(48256) := x"10e1";
    tmp(48257) := x"10e1";
    tmp(48258) := x"1101";
    tmp(48259) := x"1101";
    tmp(48260) := x"10e1";
    tmp(48261) := x"1101";
    tmp(48262) := x"1101";
    tmp(48263) := x"1101";
    tmp(48264) := x"1101";
    tmp(48265) := x"1101";
    tmp(48266) := x"1101";
    tmp(48267) := x"1101";
    tmp(48268) := x"1101";
    tmp(48269) := x"10e1";
    tmp(48270) := x"10e1";
    tmp(48271) := x"10e1";
    tmp(48272) := x"10e1";
    tmp(48273) := x"10c1";
    tmp(48274) := x"10c1";
    tmp(48275) := x"08a1";
    tmp(48276) := x"08a1";
    tmp(48277) := x"08a1";
    tmp(48278) := x"0881";
    tmp(48279) := x"0881";
    tmp(48280) := x"0881";
    tmp(48281) := x"0881";
    tmp(48282) := x"0861";
    tmp(48283) := x"0861";
    tmp(48284) := x"0861";
    tmp(48285) := x"0861";
    tmp(48286) := x"0861";
    tmp(48287) := x"0861";
    tmp(48288) := x"0861";
    tmp(48289) := x"0881";
    tmp(48290) := x"0881";
    tmp(48291) := x"0881";
    tmp(48292) := x"08a1";
    tmp(48293) := x"08a1";
    tmp(48294) := x"08a1";
    tmp(48295) := x"08a2";
    tmp(48296) := x"08a1";
    tmp(48297) := x"08a1";
    tmp(48298) := x"08a1";
    tmp(48299) := x"08a1";
    tmp(48300) := x"08a1";
    tmp(48301) := x"08c1";
    tmp(48302) := x"10e2";
    tmp(48303) := x"1103";
    tmp(48304) := x"1143";
    tmp(48305) := x"1164";
    tmp(48306) := x"1184";
    tmp(48307) := x"1164";
    tmp(48308) := x"1164";
    tmp(48309) := x"1164";
    tmp(48310) := x"1143";
    tmp(48311) := x"1143";
    tmp(48312) := x"1122";
    tmp(48313) := x"1122";
    tmp(48314) := x"1102";
    tmp(48315) := x"1102";
    tmp(48316) := x"10e1";
    tmp(48317) := x"10e1";
    tmp(48318) := x"10e1";
    tmp(48319) := x"08c1";
    tmp(48320) := x"08a1";
    tmp(48321) := x"08a0";
    tmp(48322) := x"08a0";
    tmp(48323) := x"08a0";
    tmp(48324) := x"08a0";
    tmp(48325) := x"08a0";
    tmp(48326) := x"08a0";
    tmp(48327) := x"08a0";
    tmp(48328) := x"08a0";
    tmp(48329) := x"08a0";
    tmp(48330) := x"08a0";
    tmp(48331) := x"08a0";
    tmp(48332) := x"08a0";
    tmp(48333) := x"08c0";
    tmp(48334) := x"08c0";
    tmp(48335) := x"08c0";
    tmp(48336) := x"0880";
    tmp(48337) := x"0000";
    tmp(48338) := x"0000";
    tmp(48339) := x"0820";
    tmp(48340) := x"08a0";
    tmp(48341) := x"10c0";
    tmp(48342) := x"10c0";
    tmp(48343) := x"10a0";
    tmp(48344) := x"10a0";
    tmp(48345) := x"10a0";
    tmp(48346) := x"10a0";
    tmp(48347) := x"1080";
    tmp(48348) := x"1080";
    tmp(48349) := x"0880";
    tmp(48350) := x"1080";
    tmp(48351) := x"1080";
    tmp(48352) := x"0840";
    tmp(48353) := x"0000";
    tmp(48354) := x"0000";
    tmp(48355) := x"0820";
    tmp(48356) := x"0841";
    tmp(48357) := x"0000";
    tmp(48358) := x"0000";
    tmp(48359) := x"0000";
    tmp(48360) := x"0000";
    tmp(48361) := x"0000";
    tmp(48362) := x"0000";
    tmp(48363) := x"0000";
    tmp(48364) := x"0000";
    tmp(48365) := x"0000";
    tmp(48366) := x"0000";
    tmp(48367) := x"0000";
    tmp(48368) := x"0000";
    tmp(48369) := x"0000";
    tmp(48370) := x"0000";
    tmp(48371) := x"0000";
    tmp(48372) := x"0000";
    tmp(48373) := x"0000";
    tmp(48374) := x"0000";
    tmp(48375) := x"0000";
    tmp(48376) := x"0000";
    tmp(48377) := x"0000";
    tmp(48378) := x"0000";
    tmp(48379) := x"0000";
    tmp(48380) := x"0000";
    tmp(48381) := x"0000";
    tmp(48382) := x"0000";
    tmp(48383) := x"0000";
    tmp(48384) := x"30e3";
    tmp(48385) := x"e450";
    tmp(48386) := x"eb8f";
    tmp(48387) := x"6082";
    tmp(48388) := x"3020";
    tmp(48389) := x"6882";
    tmp(48390) := x"4041";
    tmp(48391) := x"4061";
    tmp(48392) := x"4882";
    tmp(48393) := x"ba6b";
    tmp(48394) := x"8146";
    tmp(48395) := x"4042";
    tmp(48396) := x"e2ac";
    tmp(48397) := x"9987";
    tmp(48398) := x"60c4";
    tmp(48399) := x"68e4";
    tmp(48400) := x"8145";
    tmp(48401) := x"9125";
    tmp(48402) := x"a125";
    tmp(48403) := x"5841";
    tmp(48404) := x"7062";
    tmp(48405) := x"3800";
    tmp(48406) := x"5020";
    tmp(48407) := x"2800";
    tmp(48408) := x"2800";
    tmp(48409) := x"3000";
    tmp(48410) := x"3800";
    tmp(48411) := x"5000";
    tmp(48412) := x"6800";
    tmp(48413) := x"7800";
    tmp(48414) := x"7800";
    tmp(48415) := x"8800";
    tmp(48416) := x"9820";
    tmp(48417) := x"b820";
    tmp(48418) := x"c020";
    tmp(48419) := x"c020";
    tmp(48420) := x"b000";
    tmp(48421) := x"c820";
    tmp(48422) := x"c000";
    tmp(48423) := x"e020";
    tmp(48424) := x"f840";
    tmp(48425) := x"e820";
    tmp(48426) := x"d020";
    tmp(48427) := x"c040";
    tmp(48428) := x"6861";
    tmp(48429) := x"1840";
    tmp(48430) := x"1040";
    tmp(48431) := x"1040";
    tmp(48432) := x"0840";
    tmp(48433) := x"1040";
    tmp(48434) := x"0840";
    tmp(48435) := x"0840";
    tmp(48436) := x"0840";
    tmp(48437) := x"001f";
    tmp(48438) := x"001f";
    tmp(48439) := x"001f";
    tmp(48440) := x"001f";
    tmp(48441) := x"001f";
    tmp(48442) := x"001f";
    tmp(48443) := x"001f";
    tmp(48444) := x"001f";
    tmp(48445) := x"001f";
    tmp(48446) := x"001f";
    tmp(48447) := x"001f";
    tmp(48448) := x"001f";
    tmp(48449) := x"001f";
    tmp(48450) := x"001f";
    tmp(48451) := x"001f";
    tmp(48452) := x"001f";
    tmp(48453) := x"001f";
    tmp(48454) := x"001f";
    tmp(48455) := x"001f";
    tmp(48456) := x"001f";
    tmp(48457) := x"001f";
    tmp(48458) := x"001f";
    tmp(48459) := x"001f";
    tmp(48460) := x"001f";
    tmp(48461) := x"001f";
    tmp(48462) := x"001f";
    tmp(48463) := x"001f";
    tmp(48464) := x"001f";
    tmp(48465) := x"001f";
    tmp(48466) := x"001f";
    tmp(48467) := x"001f";
    tmp(48468) := x"001f";
    tmp(48469) := x"001f";
    tmp(48470) := x"001f";
    tmp(48471) := x"001f";
    tmp(48472) := x"001f";
    tmp(48473) := x"001f";
    tmp(48474) := x"001f";
    tmp(48475) := x"001f";
    tmp(48476) := x"001f";
    tmp(48477) := x"0840";
    tmp(48478) := x"0840";
    tmp(48479) := x"0840";
    tmp(48480) := x"0020";
    tmp(48481) := x"08c1";
    tmp(48482) := x"08c1";
    tmp(48483) := x"08e1";
    tmp(48484) := x"08e1";
    tmp(48485) := x"08e1";
    tmp(48486) := x"08e1";
    tmp(48487) := x"08e1";
    tmp(48488) := x"08e1";
    tmp(48489) := x"08e1";
    tmp(48490) := x"08e1";
    tmp(48491) := x"08e1";
    tmp(48492) := x"08e1";
    tmp(48493) := x"08e1";
    tmp(48494) := x"08e1";
    tmp(48495) := x"08e1";
    tmp(48496) := x"10e1";
    tmp(48497) := x"10e1";
    tmp(48498) := x"10e1";
    tmp(48499) := x"1101";
    tmp(48500) := x"10e1";
    tmp(48501) := x"1101";
    tmp(48502) := x"1101";
    tmp(48503) := x"1101";
    tmp(48504) := x"1121";
    tmp(48505) := x"1101";
    tmp(48506) := x"1121";
    tmp(48507) := x"1101";
    tmp(48508) := x"1101";
    tmp(48509) := x"1101";
    tmp(48510) := x"1101";
    tmp(48511) := x"1101";
    tmp(48512) := x"10e1";
    tmp(48513) := x"10e1";
    tmp(48514) := x"10c1";
    tmp(48515) := x"08c1";
    tmp(48516) := x"08a1";
    tmp(48517) := x"08a1";
    tmp(48518) := x"08a1";
    tmp(48519) := x"08a1";
    tmp(48520) := x"08a1";
    tmp(48521) := x"08a1";
    tmp(48522) := x"08a1";
    tmp(48523) := x"08a1";
    tmp(48524) := x"08a2";
    tmp(48525) := x"08a2";
    tmp(48526) := x"10e3";
    tmp(48527) := x"10e3";
    tmp(48528) := x"1104";
    tmp(48529) := x"1124";
    tmp(48530) := x"1125";
    tmp(48531) := x"1125";
    tmp(48532) := x"1125";
    tmp(48533) := x"1145";
    tmp(48534) := x"1145";
    tmp(48535) := x"1145";
    tmp(48536) := x"1125";
    tmp(48537) := x"1145";
    tmp(48538) := x"1145";
    tmp(48539) := x"0924";
    tmp(48540) := x"0904";
    tmp(48541) := x"0904";
    tmp(48542) := x"0925";
    tmp(48543) := x"0946";
    tmp(48544) := x"1187";
    tmp(48545) := x"0966";
    tmp(48546) := x"0945";
    tmp(48547) := x"0925";
    tmp(48548) := x"0904";
    tmp(48549) := x"08e3";
    tmp(48550) := x"08e3";
    tmp(48551) := x"0903";
    tmp(48552) := x"0923";
    tmp(48553) := x"0923";
    tmp(48554) := x"0923";
    tmp(48555) := x"1123";
    tmp(48556) := x"1144";
    tmp(48557) := x"1164";
    tmp(48558) := x"1984";
    tmp(48559) := x"19a4";
    tmp(48560) := x"1963";
    tmp(48561) := x"1143";
    tmp(48562) := x"1102";
    tmp(48563) := x"08e1";
    tmp(48564) := x"08c1";
    tmp(48565) := x"08a0";
    tmp(48566) := x"08a0";
    tmp(48567) := x"08a0";
    tmp(48568) := x"0880";
    tmp(48569) := x"0880";
    tmp(48570) := x"08a0";
    tmp(48571) := x"08a0";
    tmp(48572) := x"08a0";
    tmp(48573) := x"08a0";
    tmp(48574) := x"08a0";
    tmp(48575) := x"08c0";
    tmp(48576) := x"0840";
    tmp(48577) := x"0000";
    tmp(48578) := x"0000";
    tmp(48579) := x"0880";
    tmp(48580) := x"10a0";
    tmp(48581) := x"10a0";
    tmp(48582) := x"10a0";
    tmp(48583) := x"10a0";
    tmp(48584) := x"10a0";
    tmp(48585) := x"10a0";
    tmp(48586) := x"1080";
    tmp(48587) := x"1080";
    tmp(48588) := x"1080";
    tmp(48589) := x"0880";
    tmp(48590) := x"1080";
    tmp(48591) := x"1080";
    tmp(48592) := x"0820";
    tmp(48593) := x"0000";
    tmp(48594) := x"0000";
    tmp(48595) := x"0020";
    tmp(48596) := x"0841";
    tmp(48597) := x"0020";
    tmp(48598) := x"0000";
    tmp(48599) := x"0000";
    tmp(48600) := x"0000";
    tmp(48601) := x"0000";
    tmp(48602) := x"0000";
    tmp(48603) := x"0000";
    tmp(48604) := x"0000";
    tmp(48605) := x"0000";
    tmp(48606) := x"0000";
    tmp(48607) := x"0020";
    tmp(48608) := x"0821";
    tmp(48609) := x"0021";
    tmp(48610) := x"0000";
    tmp(48611) := x"0000";
    tmp(48612) := x"0000";
    tmp(48613) := x"0000";
    tmp(48614) := x"0000";
    tmp(48615) := x"0000";
    tmp(48616) := x"0000";
    tmp(48617) := x"0000";
    tmp(48618) := x"0000";
    tmp(48619) := x"0020";
    tmp(48620) := x"0020";
    tmp(48621) := x"0020";
    tmp(48622) := x"0000";
    tmp(48623) := x"1041";
    tmp(48624) := x"aaec";
    tmp(48625) := x"fcd5";
    tmp(48626) := x"70c4";
    tmp(48627) := x"2820";
    tmp(48628) := x"9125";
    tmp(48629) := x"4062";
    tmp(48630) := x"8966";
    tmp(48631) := x"58c3";
    tmp(48632) := x"7925";
    tmp(48633) := x"50a3";
    tmp(48634) := x"9987";
    tmp(48635) := x"a9e9";
    tmp(48636) := x"68c4";
    tmp(48637) := x"3821";
    tmp(48638) := x"5062";
    tmp(48639) := x"b1e9";
    tmp(48640) := x"b24a";
    tmp(48641) := x"3841";
    tmp(48642) := x"60a2";
    tmp(48643) := x"c9e7";
    tmp(48644) := x"6041";
    tmp(48645) := x"5020";
    tmp(48646) := x"4000";
    tmp(48647) := x"3000";
    tmp(48648) := x"3000";
    tmp(48649) := x"3000";
    tmp(48650) := x"3800";
    tmp(48651) := x"4800";
    tmp(48652) := x"6800";
    tmp(48653) := x"7800";
    tmp(48654) := x"7800";
    tmp(48655) := x"8000";
    tmp(48656) := x"a020";
    tmp(48657) := x"b820";
    tmp(48658) := x"e820";
    tmp(48659) := x"c020";
    tmp(48660) := x"a800";
    tmp(48661) := x"b800";
    tmp(48662) := x"c820";
    tmp(48663) := x"d820";
    tmp(48664) := x"f840";
    tmp(48665) := x"e840";
    tmp(48666) := x"d020";
    tmp(48667) := x"c840";
    tmp(48668) := x"7061";
    tmp(48669) := x"1840";
    tmp(48670) := x"1040";
    tmp(48671) := x"0840";
    tmp(48672) := x"0840";
    tmp(48673) := x"0840";
    tmp(48674) := x"0840";
    tmp(48675) := x"1040";
    tmp(48676) := x"0840";
    tmp(48677) := x"001f";
    tmp(48678) := x"001f";
    tmp(48679) := x"001f";
    tmp(48680) := x"001f";
    tmp(48681) := x"001f";
    tmp(48682) := x"001f";
    tmp(48683) := x"001f";
    tmp(48684) := x"001f";
    tmp(48685) := x"001f";
    tmp(48686) := x"001f";
    tmp(48687) := x"001f";
    tmp(48688) := x"001f";
    tmp(48689) := x"001f";
    tmp(48690) := x"001f";
    tmp(48691) := x"001f";
    tmp(48692) := x"001f";
    tmp(48693) := x"001f";
    tmp(48694) := x"001f";
    tmp(48695) := x"001f";
    tmp(48696) := x"001f";
    tmp(48697) := x"001f";
    tmp(48698) := x"001f";
    tmp(48699) := x"001f";
    tmp(48700) := x"001f";
    tmp(48701) := x"001f";
    tmp(48702) := x"001f";
    tmp(48703) := x"001f";
    tmp(48704) := x"001f";
    tmp(48705) := x"001f";
    tmp(48706) := x"001f";
    tmp(48707) := x"001f";
    tmp(48708) := x"001f";
    tmp(48709) := x"001f";
    tmp(48710) := x"001f";
    tmp(48711) := x"001f";
    tmp(48712) := x"001f";
    tmp(48713) := x"001f";
    tmp(48714) := x"001f";
    tmp(48715) := x"001f";
    tmp(48716) := x"001f";
    tmp(48717) := x"0840";
    tmp(48718) := x"0840";
    tmp(48719) := x"0840";
    tmp(48720) := x"0020";
    tmp(48721) := x"08c1";
    tmp(48722) := x"08c1";
    tmp(48723) := x"08e1";
    tmp(48724) := x"08e1";
    tmp(48725) := x"08e1";
    tmp(48726) := x"08e1";
    tmp(48727) := x"08e1";
    tmp(48728) := x"08e1";
    tmp(48729) := x"08e1";
    tmp(48730) := x"08e1";
    tmp(48731) := x"08e1";
    tmp(48732) := x"08c1";
    tmp(48733) := x"08e1";
    tmp(48734) := x"08e1";
    tmp(48735) := x"08c1";
    tmp(48736) := x"08c1";
    tmp(48737) := x"08e1";
    tmp(48738) := x"08e1";
    tmp(48739) := x"10e1";
    tmp(48740) := x"10e1";
    tmp(48741) := x"1101";
    tmp(48742) := x"1101";
    tmp(48743) := x"1121";
    tmp(48744) := x"1101";
    tmp(48745) := x"1121";
    tmp(48746) := x"1121";
    tmp(48747) := x"1101";
    tmp(48748) := x"1101";
    tmp(48749) := x"1101";
    tmp(48750) := x"1101";
    tmp(48751) := x"1101";
    tmp(48752) := x"10e1";
    tmp(48753) := x"10e1";
    tmp(48754) := x"08e1";
    tmp(48755) := x"08e2";
    tmp(48756) := x"08e2";
    tmp(48757) := x"0902";
    tmp(48758) := x"1103";
    tmp(48759) := x"1124";
    tmp(48760) := x"1145";
    tmp(48761) := x"1145";
    tmp(48762) := x"1104";
    tmp(48763) := x"08c3";
    tmp(48764) := x"08a2";
    tmp(48765) := x"0882";
    tmp(48766) := x"0882";
    tmp(48767) := x"0861";
    tmp(48768) := x"0861";
    tmp(48769) := x"0041";
    tmp(48770) := x"0041";
    tmp(48771) := x"0041";
    tmp(48772) := x"0041";
    tmp(48773) := x"0041";
    tmp(48774) := x"0041";
    tmp(48775) := x"0041";
    tmp(48776) := x"0041";
    tmp(48777) := x"0061";
    tmp(48778) := x"0061";
    tmp(48779) := x"0082";
    tmp(48780) := x"0082";
    tmp(48781) := x"08a2";
    tmp(48782) := x"08a3";
    tmp(48783) := x"08c3";
    tmp(48784) := x"08e4";
    tmp(48785) := x"08e4";
    tmp(48786) := x"0905";
    tmp(48787) := x"08e4";
    tmp(48788) := x"08a3";
    tmp(48789) := x"08a2";
    tmp(48790) := x"0882";
    tmp(48791) := x"0881";
    tmp(48792) := x"0881";
    tmp(48793) := x"0060";
    tmp(48794) := x"0060";
    tmp(48795) := x"0060";
    tmp(48796) := x"0040";
    tmp(48797) := x"0040";
    tmp(48798) := x"0040";
    tmp(48799) := x"0060";
    tmp(48800) := x"0861";
    tmp(48801) := x"08a1";
    tmp(48802) := x"08c2";
    tmp(48803) := x"1102";
    tmp(48804) := x"1123";
    tmp(48805) := x"1102";
    tmp(48806) := x"10e2";
    tmp(48807) := x"10c1";
    tmp(48808) := x"08a1";
    tmp(48809) := x"08a0";
    tmp(48810) := x"08a0";
    tmp(48811) := x"08a0";
    tmp(48812) := x"0880";
    tmp(48813) := x"08a0";
    tmp(48814) := x"08a0";
    tmp(48815) := x"08a0";
    tmp(48816) := x"0020";
    tmp(48817) := x"0000";
    tmp(48818) := x"0840";
    tmp(48819) := x"10a0";
    tmp(48820) := x"08a0";
    tmp(48821) := x"10a0";
    tmp(48822) := x"10a0";
    tmp(48823) := x"10a0";
    tmp(48824) := x"1080";
    tmp(48825) := x"1080";
    tmp(48826) := x"1080";
    tmp(48827) := x"1080";
    tmp(48828) := x"1080";
    tmp(48829) := x"1080";
    tmp(48830) := x"1080";
    tmp(48831) := x"1080";
    tmp(48832) := x"0820";
    tmp(48833) := x"0000";
    tmp(48834) := x"0000";
    tmp(48835) := x"0020";
    tmp(48836) := x"0020";
    tmp(48837) := x"0841";
    tmp(48838) := x"0020";
    tmp(48839) := x"0000";
    tmp(48840) := x"0000";
    tmp(48841) := x"0000";
    tmp(48842) := x"0000";
    tmp(48843) := x"0000";
    tmp(48844) := x"0000";
    tmp(48845) := x"0000";
    tmp(48846) := x"0000";
    tmp(48847) := x"0020";
    tmp(48848) := x"0021";
    tmp(48849) := x"0000";
    tmp(48850) := x"0000";
    tmp(48851) := x"0000";
    tmp(48852) := x"0000";
    tmp(48853) := x"0000";
    tmp(48854) := x"0000";
    tmp(48855) := x"0000";
    tmp(48856) := x"0000";
    tmp(48857) := x"0000";
    tmp(48858) := x"0000";
    tmp(48859) := x"0000";
    tmp(48860) := x"0000";
    tmp(48861) := x"0020";
    tmp(48862) := x"0820";
    tmp(48863) := x"38e3";
    tmp(48864) := x"e472";
    tmp(48865) := x"91a7";
    tmp(48866) := x"3020";
    tmp(48867) := x"9945";
    tmp(48868) := x"b1e8";
    tmp(48869) := x"6104";
    tmp(48870) := x"7946";
    tmp(48871) := x"4882";
    tmp(48872) := x"8166";
    tmp(48873) := x"4041";
    tmp(48874) := x"4862";
    tmp(48875) := x"7925";
    tmp(48876) := x"4041";
    tmp(48877) := x"80e4";
    tmp(48878) := x"b1c7";
    tmp(48879) := x"9187";
    tmp(48880) := x"9187";
    tmp(48881) := x"cacc";
    tmp(48882) := x"60a2";
    tmp(48883) := x"8904";
    tmp(48884) := x"9125";
    tmp(48885) := x"3820";
    tmp(48886) := x"98a2";
    tmp(48887) := x"3000";
    tmp(48888) := x"3800";
    tmp(48889) := x"4000";
    tmp(48890) := x"4000";
    tmp(48891) := x"5000";
    tmp(48892) := x"6800";
    tmp(48893) := x"7800";
    tmp(48894) := x"7800";
    tmp(48895) := x"9000";
    tmp(48896) := x"a820";
    tmp(48897) := x"c020";
    tmp(48898) := x"e020";
    tmp(48899) := x"c020";
    tmp(48900) := x"a800";
    tmp(48901) := x"b800";
    tmp(48902) := x"b800";
    tmp(48903) := x"c820";
    tmp(48904) := x"e820";
    tmp(48905) := x"e820";
    tmp(48906) := x"d820";
    tmp(48907) := x"d040";
    tmp(48908) := x"6861";
    tmp(48909) := x"1840";
    tmp(48910) := x"1040";
    tmp(48911) := x"1040";
    tmp(48912) := x"0840";
    tmp(48913) := x"0840";
    tmp(48914) := x"0840";
    tmp(48915) := x"0840";
    tmp(48916) := x"0840";
    tmp(48917) := x"001f";
    tmp(48918) := x"001f";
    tmp(48919) := x"001f";
    tmp(48920) := x"001f";
    tmp(48921) := x"001f";
    tmp(48922) := x"001f";
    tmp(48923) := x"001f";
    tmp(48924) := x"001f";
    tmp(48925) := x"001f";
    tmp(48926) := x"001f";
    tmp(48927) := x"001f";
    tmp(48928) := x"001f";
    tmp(48929) := x"001f";
    tmp(48930) := x"001f";
    tmp(48931) := x"001f";
    tmp(48932) := x"001f";
    tmp(48933) := x"001f";
    tmp(48934) := x"001f";
    tmp(48935) := x"001f";
    tmp(48936) := x"001f";
    tmp(48937) := x"001f";
    tmp(48938) := x"001f";
    tmp(48939) := x"001f";
    tmp(48940) := x"001f";
    tmp(48941) := x"001f";
    tmp(48942) := x"001f";
    tmp(48943) := x"001f";
    tmp(48944) := x"001f";
    tmp(48945) := x"001f";
    tmp(48946) := x"001f";
    tmp(48947) := x"001f";
    tmp(48948) := x"001f";
    tmp(48949) := x"001f";
    tmp(48950) := x"001f";
    tmp(48951) := x"001f";
    tmp(48952) := x"001f";
    tmp(48953) := x"001f";
    tmp(48954) := x"001f";
    tmp(48955) := x"001f";
    tmp(48956) := x"001f";
    tmp(48957) := x"0840";
    tmp(48958) := x"0840";
    tmp(48959) := x"0840";
    tmp(48960) := x"0000";
    tmp(48961) := x"08c1";
    tmp(48962) := x"08c1";
    tmp(48963) := x"08e1";
    tmp(48964) := x"08e1";
    tmp(48965) := x"08e1";
    tmp(48966) := x"08e1";
    tmp(48967) := x"08e1";
    tmp(48968) := x"08e1";
    tmp(48969) := x"08e1";
    tmp(48970) := x"08e1";
    tmp(48971) := x"08e1";
    tmp(48972) := x"08e1";
    tmp(48973) := x"08e1";
    tmp(48974) := x"08e1";
    tmp(48975) := x"08e1";
    tmp(48976) := x"08e1";
    tmp(48977) := x"08e1";
    tmp(48978) := x"08e1";
    tmp(48979) := x"08e1";
    tmp(48980) := x"10e1";
    tmp(48981) := x"10e1";
    tmp(48982) := x"1101";
    tmp(48983) := x"1101";
    tmp(48984) := x"1101";
    tmp(48985) := x"1101";
    tmp(48986) := x"1121";
    tmp(48987) := x"1121";
    tmp(48988) := x"1121";
    tmp(48989) := x"1121";
    tmp(48990) := x"1122";
    tmp(48991) := x"1122";
    tmp(48992) := x"1123";
    tmp(48993) := x"0923";
    tmp(48994) := x"1144";
    tmp(48995) := x"0945";
    tmp(48996) := x"0945";
    tmp(48997) := x"0925";
    tmp(48998) := x"08e4";
    tmp(48999) := x"08a2";
    tmp(49000) := x"0061";
    tmp(49001) := x"0041";
    tmp(49002) := x"0021";
    tmp(49003) := x"0020";
    tmp(49004) := x"0020";
    tmp(49005) := x"0020";
    tmp(49006) := x"0020";
    tmp(49007) := x"0021";
    tmp(49008) := x"0041";
    tmp(49009) := x"0041";
    tmp(49010) := x"0041";
    tmp(49011) := x"0041";
    tmp(49012) := x"0041";
    tmp(49013) := x"0021";
    tmp(49014) := x"0021";
    tmp(49015) := x"0021";
    tmp(49016) := x"0021";
    tmp(49017) := x"0041";
    tmp(49018) := x"0041";
    tmp(49019) := x"0021";
    tmp(49020) := x"0041";
    tmp(49021) := x"0041";
    tmp(49022) := x"0041";
    tmp(49023) := x"0061";
    tmp(49024) := x"0061";
    tmp(49025) := x"0061";
    tmp(49026) := x"0062";
    tmp(49027) := x"0082";
    tmp(49028) := x"0082";
    tmp(49029) := x"00a2";
    tmp(49030) := x"08a3";
    tmp(49031) := x"08a2";
    tmp(49032) := x"08c2";
    tmp(49033) := x"08c2";
    tmp(49034) := x"08e1";
    tmp(49035) := x"08e1";
    tmp(49036) := x"10e1";
    tmp(49037) := x"10e1";
    tmp(49038) := x"10c1";
    tmp(49039) := x"08a1";
    tmp(49040) := x"08a0";
    tmp(49041) := x"0880";
    tmp(49042) := x"0860";
    tmp(49043) := x"0860";
    tmp(49044) := x"0860";
    tmp(49045) := x"0881";
    tmp(49046) := x"08a1";
    tmp(49047) := x"10c1";
    tmp(49048) := x"18e1";
    tmp(49049) := x"10a1";
    tmp(49050) := x"10a0";
    tmp(49051) := x"10a0";
    tmp(49052) := x"10a0";
    tmp(49053) := x"1080";
    tmp(49054) := x"10a0";
    tmp(49055) := x"0880";
    tmp(49056) := x"0020";
    tmp(49057) := x"0020";
    tmp(49058) := x"1080";
    tmp(49059) := x"0880";
    tmp(49060) := x"0880";
    tmp(49061) := x"0880";
    tmp(49062) := x"1080";
    tmp(49063) := x"1080";
    tmp(49064) := x"1080";
    tmp(49065) := x"1080";
    tmp(49066) := x"1080";
    tmp(49067) := x"0880";
    tmp(49068) := x"1080";
    tmp(49069) := x"1080";
    tmp(49070) := x"1060";
    tmp(49071) := x"1060";
    tmp(49072) := x"0820";
    tmp(49073) := x"0000";
    tmp(49074) := x"0000";
    tmp(49075) := x"0000";
    tmp(49076) := x"0000";
    tmp(49077) := x"0020";
    tmp(49078) := x"0020";
    tmp(49079) := x"0020";
    tmp(49080) := x"0020";
    tmp(49081) := x"0000";
    tmp(49082) := x"0020";
    tmp(49083) := x"0000";
    tmp(49084) := x"0000";
    tmp(49085) := x"0000";
    tmp(49086) := x"0000";
    tmp(49087) := x"0000";
    tmp(49088) := x"0000";
    tmp(49089) := x"0000";
    tmp(49090) := x"0000";
    tmp(49091) := x"0000";
    tmp(49092) := x"0000";
    tmp(49093) := x"0000";
    tmp(49094) := x"0000";
    tmp(49095) := x"0000";
    tmp(49096) := x"0000";
    tmp(49097) := x"0000";
    tmp(49098) := x"0000";
    tmp(49099) := x"0000";
    tmp(49100) := x"0000";
    tmp(49101) := x"0000";
    tmp(49102) := x"1020";
    tmp(49103) := x"5124";
    tmp(49104) := x"9186";
    tmp(49105) := x"3821";
    tmp(49106) := x"4041";
    tmp(49107) := x"dacc";
    tmp(49108) := x"3862";
    tmp(49109) := x"8186";
    tmp(49110) := x"6904";
    tmp(49111) := x"4061";
    tmp(49112) := x"daec";
    tmp(49113) := x"a1c8";
    tmp(49114) := x"5882";
    tmp(49115) := x"c1e8";
    tmp(49116) := x"f34e";
    tmp(49117) := x"8125";
    tmp(49118) := x"2820";
    tmp(49119) := x"2800";
    tmp(49120) := x"2820";
    tmp(49121) := x"3841";
    tmp(49122) := x"3841";
    tmp(49123) := x"2820";
    tmp(49124) := x"78c3";
    tmp(49125) := x"5041";
    tmp(49126) := x"4821";
    tmp(49127) := x"3000";
    tmp(49128) := x"3000";
    tmp(49129) := x"4000";
    tmp(49130) := x"4000";
    tmp(49131) := x"5000";
    tmp(49132) := x"6000";
    tmp(49133) := x"7800";
    tmp(49134) := x"8800";
    tmp(49135) := x"9800";
    tmp(49136) := x"a020";
    tmp(49137) := x"c820";
    tmp(49138) := x"f020";
    tmp(49139) := x"c820";
    tmp(49140) := x"a800";
    tmp(49141) := x"c020";
    tmp(49142) := x"c020";
    tmp(49143) := x"d020";
    tmp(49144) := x"e020";
    tmp(49145) := x"e020";
    tmp(49146) := x"e820";
    tmp(49147) := x"d040";
    tmp(49148) := x"5860";
    tmp(49149) := x"1840";
    tmp(49150) := x"1040";
    tmp(49151) := x"0840";
    tmp(49152) := x"0840";
    tmp(49153) := x"0840";
    tmp(49154) := x"0840";
    tmp(49155) := x"0840";
    tmp(49156) := x"0840";
    tmp(49157) := x"0840";
    tmp(49158) := x"0840";
    tmp(49159) := x"0840";
    tmp(49160) := x"0840";
    tmp(49161) := x"0840";
    tmp(49162) := x"0840";
    tmp(49163) := x"0840";
    tmp(49164) := x"0840";
    tmp(49165) := x"0840";
    tmp(49166) := x"0840";
    tmp(49167) := x"0840";
    tmp(49168) := x"0840";
    tmp(49169) := x"0840";
    tmp(49170) := x"0840";
    tmp(49171) := x"0840";
    tmp(49172) := x"0840";
    tmp(49173) := x"0840";
    tmp(49174) := x"0840";
    tmp(49175) := x"0840";
    tmp(49176) := x"0840";
    tmp(49177) := x"0840";
    tmp(49178) := x"0840";
    tmp(49179) := x"0840";
    tmp(49180) := x"0840";
    tmp(49181) := x"0840";
    tmp(49182) := x"0840";
    tmp(49183) := x"0840";
    tmp(49184) := x"0840";
    tmp(49185) := x"0840";
    tmp(49186) := x"0840";
    tmp(49187) := x"0840";
    tmp(49188) := x"0840";
    tmp(49189) := x"0840";
    tmp(49190) := x"0840";
    tmp(49191) := x"0840";
    tmp(49192) := x"0840";
    tmp(49193) := x"0840";
    tmp(49194) := x"0840";
    tmp(49195) := x"0840";
    tmp(49196) := x"0840";
    tmp(49197) := x"0840";
    tmp(49198) := x"0840";
    tmp(49199) := x"0840";
    tmp(49200) := x"0000";
    tmp(49201) := x"08c1";
    tmp(49202) := x"08c1";
    tmp(49203) := x"08e1";
    tmp(49204) := x"08e1";
    tmp(49205) := x"08e1";
    tmp(49206) := x"08c1";
    tmp(49207) := x"08c0";
    tmp(49208) := x"08e1";
    tmp(49209) := x"08e1";
    tmp(49210) := x"08e1";
    tmp(49211) := x"08e1";
    tmp(49212) := x"08e1";
    tmp(49213) := x"1101";
    tmp(49214) := x"1101";
    tmp(49215) := x"10e1";
    tmp(49216) := x"08e1";
    tmp(49217) := x"08e1";
    tmp(49218) := x"08e1";
    tmp(49219) := x"08e1";
    tmp(49220) := x"10e1";
    tmp(49221) := x"10e1";
    tmp(49222) := x"1101";
    tmp(49223) := x"10e1";
    tmp(49224) := x"1101";
    tmp(49225) := x"1101";
    tmp(49226) := x"1121";
    tmp(49227) := x"1122";
    tmp(49228) := x"1122";
    tmp(49229) := x"1143";
    tmp(49230) := x"0944";
    tmp(49231) := x"0965";
    tmp(49232) := x"0966";
    tmp(49233) := x"0925";
    tmp(49234) := x"08c3";
    tmp(49235) := x"0082";
    tmp(49236) := x"0041";
    tmp(49237) := x"0020";
    tmp(49238) := x"0020";
    tmp(49239) := x"0020";
    tmp(49240) := x"0021";
    tmp(49241) := x"0041";
    tmp(49242) := x"0041";
    tmp(49243) := x"0041";
    tmp(49244) := x"0061";
    tmp(49245) := x"0082";
    tmp(49246) := x"0083";
    tmp(49247) := x"00a3";
    tmp(49248) := x"08c4";
    tmp(49249) := x"08c4";
    tmp(49250) := x"08e5";
    tmp(49251) := x"08e5";
    tmp(49252) := x"08e5";
    tmp(49253) := x"08e5";
    tmp(49254) := x"0906";
    tmp(49255) := x"0906";
    tmp(49256) := x"0906";
    tmp(49257) := x"0926";
    tmp(49258) := x"0926";
    tmp(49259) := x"0926";
    tmp(49260) := x"0906";
    tmp(49261) := x"0906";
    tmp(49262) := x"0906";
    tmp(49263) := x"0905";
    tmp(49264) := x"0905";
    tmp(49265) := x"08e5";
    tmp(49266) := x"08c4";
    tmp(49267) := x"08c3";
    tmp(49268) := x"08c3";
    tmp(49269) := x"08a3";
    tmp(49270) := x"0082";
    tmp(49271) := x"0082";
    tmp(49272) := x"0062";
    tmp(49273) := x"0061";
    tmp(49274) := x"0041";
    tmp(49275) := x"0040";
    tmp(49276) := x"0860";
    tmp(49277) := x"0880";
    tmp(49278) := x"10a0";
    tmp(49279) := x"10c0";
    tmp(49280) := x"10e1";
    tmp(49281) := x"18c1";
    tmp(49282) := x"18c1";
    tmp(49283) := x"18c1";
    tmp(49284) := x"18c1";
    tmp(49285) := x"18e1";
    tmp(49286) := x"18a1";
    tmp(49287) := x"1061";
    tmp(49288) := x"1060";
    tmp(49289) := x"1060";
    tmp(49290) := x"1060";
    tmp(49291) := x"1880";
    tmp(49292) := x"20c0";
    tmp(49293) := x"20c0";
    tmp(49294) := x"20c0";
    tmp(49295) := x"1060";
    tmp(49296) := x"0840";
    tmp(49297) := x"1080";
    tmp(49298) := x"1080";
    tmp(49299) := x"1080";
    tmp(49300) := x"0880";
    tmp(49301) := x"1080";
    tmp(49302) := x"1080";
    tmp(49303) := x"1080";
    tmp(49304) := x"1080";
    tmp(49305) := x"1080";
    tmp(49306) := x"1080";
    tmp(49307) := x"1080";
    tmp(49308) := x"1060";
    tmp(49309) := x"1060";
    tmp(49310) := x"0860";
    tmp(49311) := x"0860";
    tmp(49312) := x"0020";
    tmp(49313) := x"0000";
    tmp(49314) := x"0000";
    tmp(49315) := x"0000";
    tmp(49316) := x"0000";
    tmp(49317) := x"0000";
    tmp(49318) := x"0000";
    tmp(49319) := x"0000";
    tmp(49320) := x"0000";
    tmp(49321) := x"0000";
    tmp(49322) := x"0000";
    tmp(49323) := x"0000";
    tmp(49324) := x"0820";
    tmp(49325) := x"0841";
    tmp(49326) := x"0820";
    tmp(49327) := x"0821";
    tmp(49328) := x"0020";
    tmp(49329) := x"0000";
    tmp(49330) := x"0000";
    tmp(49331) := x"0000";
    tmp(49332) := x"0000";
    tmp(49333) := x"0000";
    tmp(49334) := x"0020";
    tmp(49335) := x"0020";
    tmp(49336) := x"0000";
    tmp(49337) := x"0000";
    tmp(49338) := x"0000";
    tmp(49339) := x"0000";
    tmp(49340) := x"1041";
    tmp(49341) := x"1861";
    tmp(49342) := x"38a2";
    tmp(49343) := x"60a3";
    tmp(49344) := x"3020";
    tmp(49345) := x"3821";
    tmp(49346) := x"ba49";
    tmp(49347) := x"8166";
    tmp(49348) := x"8966";
    tmp(49349) := x"ba4a";
    tmp(49350) := x"60c3";
    tmp(49351) := x"68c3";
    tmp(49352) := x"60e4";
    tmp(49353) := x"c2ac";
    tmp(49354) := x"a9e8";
    tmp(49355) := x"3841";
    tmp(49356) := x"3021";
    tmp(49357) := x"3021";
    tmp(49358) := x"2800";
    tmp(49359) := x"4021";
    tmp(49360) := x"88e3";
    tmp(49361) := x"8904";
    tmp(49362) := x"70c3";
    tmp(49363) := x"c208";
    tmp(49364) := x"70c3";
    tmp(49365) := x"3841";
    tmp(49366) := x"3020";
    tmp(49367) := x"3820";
    tmp(49368) := x"3000";
    tmp(49369) := x"4000";
    tmp(49370) := x"4800";
    tmp(49371) := x"5800";
    tmp(49372) := x"6000";
    tmp(49373) := x"7820";
    tmp(49374) := x"9820";
    tmp(49375) := x"a020";
    tmp(49376) := x"a820";
    tmp(49377) := x"c820";
    tmp(49378) := x"e020";
    tmp(49379) := x"c820";
    tmp(49380) := x"a800";
    tmp(49381) := x"c020";
    tmp(49382) := x"d020";
    tmp(49383) := x"d820";
    tmp(49384) := x"d820";
    tmp(49385) := x"d820";
    tmp(49386) := x"e820";
    tmp(49387) := x"e840";
    tmp(49388) := x"7061";
    tmp(49389) := x"1840";
    tmp(49390) := x"0840";
    tmp(49391) := x"0840";
    tmp(49392) := x"0840";
    tmp(49393) := x"0840";
    tmp(49394) := x"0840";
    tmp(49395) := x"0840";
    tmp(49396) := x"0840";
    tmp(49397) := x"0840";
    tmp(49398) := x"0840";
    tmp(49399) := x"0840";
    tmp(49400) := x"0840";
    tmp(49401) := x"0840";
    tmp(49402) := x"0840";
    tmp(49403) := x"0840";
    tmp(49404) := x"0840";
    tmp(49405) := x"0840";
    tmp(49406) := x"0840";
    tmp(49407) := x"0840";
    tmp(49408) := x"0840";
    tmp(49409) := x"0840";
    tmp(49410) := x"0840";
    tmp(49411) := x"0840";
    tmp(49412) := x"0840";
    tmp(49413) := x"0840";
    tmp(49414) := x"0840";
    tmp(49415) := x"0840";
    tmp(49416) := x"0840";
    tmp(49417) := x"0840";
    tmp(49418) := x"0840";
    tmp(49419) := x"0840";
    tmp(49420) := x"0840";
    tmp(49421) := x"0840";
    tmp(49422) := x"0840";
    tmp(49423) := x"0840";
    tmp(49424) := x"0840";
    tmp(49425) := x"0840";
    tmp(49426) := x"0840";
    tmp(49427) := x"0840";
    tmp(49428) := x"0840";
    tmp(49429) := x"0840";
    tmp(49430) := x"0840";
    tmp(49431) := x"0840";
    tmp(49432) := x"0840";
    tmp(49433) := x"0840";
    tmp(49434) := x"0840";
    tmp(49435) := x"0840";
    tmp(49436) := x"0840";
    tmp(49437) := x"0840";
    tmp(49438) := x"0840";
    tmp(49439) := x"0840";
    tmp(49440) := x"0000";
    tmp(49441) := x"08a0";
    tmp(49442) := x"08c0";
    tmp(49443) := x"08c1";
    tmp(49444) := x"08e1";
    tmp(49445) := x"08e1";
    tmp(49446) := x"08c0";
    tmp(49447) := x"08c0";
    tmp(49448) := x"08c1";
    tmp(49449) := x"08c1";
    tmp(49450) := x"08e1";
    tmp(49451) := x"08e1";
    tmp(49452) := x"10e1";
    tmp(49453) := x"1101";
    tmp(49454) := x"1101";
    tmp(49455) := x"10e1";
    tmp(49456) := x"10e1";
    tmp(49457) := x"10e1";
    tmp(49458) := x"1101";
    tmp(49459) := x"10e1";
    tmp(49460) := x"10e1";
    tmp(49461) := x"1101";
    tmp(49462) := x"1101";
    tmp(49463) := x"1101";
    tmp(49464) := x"1102";
    tmp(49465) := x"0902";
    tmp(49466) := x"0903";
    tmp(49467) := x"08e3";
    tmp(49468) := x"08e4";
    tmp(49469) := x"08e4";
    tmp(49470) := x"08a3";
    tmp(49471) := x"0082";
    tmp(49472) := x"0041";
    tmp(49473) := x"0041";
    tmp(49474) := x"0041";
    tmp(49475) := x"0041";
    tmp(49476) := x"0041";
    tmp(49477) := x"0062";
    tmp(49478) := x"0082";
    tmp(49479) := x"0082";
    tmp(49480) := x"0082";
    tmp(49481) := x"0082";
    tmp(49482) := x"0082";
    tmp(49483) := x"0082";
    tmp(49484) := x"0082";
    tmp(49485) := x"0082";
    tmp(49486) := x"0082";
    tmp(49487) := x"0082";
    tmp(49488) := x"0062";
    tmp(49489) := x"0062";
    tmp(49490) := x"0062";
    tmp(49491) := x"0082";
    tmp(49492) := x"0082";
    tmp(49493) := x"0082";
    tmp(49494) := x"0082";
    tmp(49495) := x"0082";
    tmp(49496) := x"0082";
    tmp(49497) := x"0082";
    tmp(49498) := x"0082";
    tmp(49499) := x"00a3";
    tmp(49500) := x"00a3";
    tmp(49501) := x"00a3";
    tmp(49502) := x"08a3";
    tmp(49503) := x"08c4";
    tmp(49504) := x"08e5";
    tmp(49505) := x"0905";
    tmp(49506) := x"0906";
    tmp(49507) := x"0905";
    tmp(49508) := x"1146";
    tmp(49509) := x"1167";
    tmp(49510) := x"1147";
    tmp(49511) := x"0926";
    tmp(49512) := x"0926";
    tmp(49513) := x"08e5";
    tmp(49514) := x"0862";
    tmp(49515) := x"0820";
    tmp(49516) := x"1040";
    tmp(49517) := x"0840";
    tmp(49518) := x"0840";
    tmp(49519) := x"0840";
    tmp(49520) := x"0840";
    tmp(49521) := x"0840";
    tmp(49522) := x"0840";
    tmp(49523) := x"0840";
    tmp(49524) := x"0840";
    tmp(49525) := x"1040";
    tmp(49526) := x"1061";
    tmp(49527) := x"1081";
    tmp(49528) := x"1081";
    tmp(49529) := x"1060";
    tmp(49530) := x"1840";
    tmp(49531) := x"1860";
    tmp(49532) := x"2081";
    tmp(49533) := x"28c1";
    tmp(49534) := x"28c1";
    tmp(49535) := x"20a1";
    tmp(49536) := x"28a1";
    tmp(49537) := x"28c1";
    tmp(49538) := x"20a1";
    tmp(49539) := x"1881";
    tmp(49540) := x"1060";
    tmp(49541) := x"1060";
    tmp(49542) := x"1060";
    tmp(49543) := x"1060";
    tmp(49544) := x"1060";
    tmp(49545) := x"0860";
    tmp(49546) := x"1060";
    tmp(49547) := x"1060";
    tmp(49548) := x"1060";
    tmp(49549) := x"0860";
    tmp(49550) := x"0860";
    tmp(49551) := x"0840";
    tmp(49552) := x"0020";
    tmp(49553) := x"0000";
    tmp(49554) := x"0000";
    tmp(49555) := x"0000";
    tmp(49556) := x"0000";
    tmp(49557) := x"0000";
    tmp(49558) := x"0000";
    tmp(49559) := x"0000";
    tmp(49560) := x"0000";
    tmp(49561) := x"0000";
    tmp(49562) := x"0000";
    tmp(49563) := x"0000";
    tmp(49564) := x"0000";
    tmp(49565) := x"0000";
    tmp(49566) := x"0000";
    tmp(49567) := x"0020";
    tmp(49568) := x"0841";
    tmp(49569) := x"0820";
    tmp(49570) := x"0000";
    tmp(49571) := x"0000";
    tmp(49572) := x"0000";
    tmp(49573) := x"0000";
    tmp(49574) := x"0020";
    tmp(49575) := x"0020";
    tmp(49576) := x"0000";
    tmp(49577) := x"0000";
    tmp(49578) := x"0000";
    tmp(49579) := x"1021";
    tmp(49580) := x"2081";
    tmp(49581) := x"3082";
    tmp(49582) := x"4082";
    tmp(49583) := x"4021";
    tmp(49584) := x"2800";
    tmp(49585) := x"5082";
    tmp(49586) := x"db6e";
    tmp(49587) := x"7166";
    tmp(49588) := x"b28b";
    tmp(49589) := x"aa09";
    tmp(49590) := x"58c3";
    tmp(49591) := x"8166";
    tmp(49592) := x"7125";
    tmp(49593) := x"8986";
    tmp(49594) := x"a9e8";
    tmp(49595) := x"b1a8";
    tmp(49596) := x"ca6b";
    tmp(49597) := x"ba4a";
    tmp(49598) := x"8925";
    tmp(49599) := x"68a3";
    tmp(49600) := x"3021";
    tmp(49601) := x"60a2";
    tmp(49602) := x"c249";
    tmp(49603) := x"8145";
    tmp(49604) := x"8925";
    tmp(49605) := x"70c3";
    tmp(49606) := x"2820";
    tmp(49607) := x"4020";
    tmp(49608) := x"3000";
    tmp(49609) := x"4800";
    tmp(49610) := x"5800";
    tmp(49611) := x"6000";
    tmp(49612) := x"6000";
    tmp(49613) := x"7800";
    tmp(49614) := x"9820";
    tmp(49615) := x"a820";
    tmp(49616) := x"a020";
    tmp(49617) := x"b820";
    tmp(49618) := x"d820";
    tmp(49619) := x"c820";
    tmp(49620) := x"b000";
    tmp(49621) := x"e820";
    tmp(49622) := x"d820";
    tmp(49623) := x"c820";
    tmp(49624) := x"e020";
    tmp(49625) := x"c820";
    tmp(49626) := x"e820";
    tmp(49627) := x"f841";
    tmp(49628) := x"7861";
    tmp(49629) := x"1840";
    tmp(49630) := x"0840";
    tmp(49631) := x"0840";
    tmp(49632) := x"0840";
    tmp(49633) := x"0840";
    tmp(49634) := x"0840";
    tmp(49635) := x"0840";
    tmp(49636) := x"0840";
    tmp(49637) := x"0840";
    tmp(49638) := x"0840";
    tmp(49639) := x"0840";
    tmp(49640) := x"0840";
    tmp(49641) := x"0840";
    tmp(49642) := x"0840";
    tmp(49643) := x"0840";
    tmp(49644) := x"0840";
    tmp(49645) := x"0840";
    tmp(49646) := x"0840";
    tmp(49647) := x"0840";
    tmp(49648) := x"0840";
    tmp(49649) := x"0840";
    tmp(49650) := x"0840";
    tmp(49651) := x"0840";
    tmp(49652) := x"0840";
    tmp(49653) := x"0840";
    tmp(49654) := x"0840";
    tmp(49655) := x"0840";
    tmp(49656) := x"0840";
    tmp(49657) := x"0840";
    tmp(49658) := x"0840";
    tmp(49659) := x"0840";
    tmp(49660) := x"0840";
    tmp(49661) := x"0840";
    tmp(49662) := x"0840";
    tmp(49663) := x"0840";
    tmp(49664) := x"0840";
    tmp(49665) := x"0840";
    tmp(49666) := x"0840";
    tmp(49667) := x"0840";
    tmp(49668) := x"0840";
    tmp(49669) := x"0840";
    tmp(49670) := x"0840";
    tmp(49671) := x"0840";
    tmp(49672) := x"0840";
    tmp(49673) := x"0840";
    tmp(49674) := x"0840";
    tmp(49675) := x"0840";
    tmp(49676) := x"0840";
    tmp(49677) := x"0840";
    tmp(49678) := x"0840";
    tmp(49679) := x"0840";
    tmp(49680) := x"0000";
    tmp(49681) := x"08a0";
    tmp(49682) := x"08a0";
    tmp(49683) := x"08c0";
    tmp(49684) := x"08c1";
    tmp(49685) := x"08c1";
    tmp(49686) := x"08c0";
    tmp(49687) := x"08c0";
    tmp(49688) := x"08c1";
    tmp(49689) := x"08e1";
    tmp(49690) := x"08e1";
    tmp(49691) := x"08e1";
    tmp(49692) := x"08e1";
    tmp(49693) := x"08e1";
    tmp(49694) := x"1101";
    tmp(49695) := x"10e1";
    tmp(49696) := x"1101";
    tmp(49697) := x"1101";
    tmp(49698) := x"1101";
    tmp(49699) := x"1101";
    tmp(49700) := x"1101";
    tmp(49701) := x"1102";
    tmp(49702) := x"08e2";
    tmp(49703) := x"08e2";
    tmp(49704) := x"08a2";
    tmp(49705) := x"0082";
    tmp(49706) := x"0062";
    tmp(49707) := x"0061";
    tmp(49708) := x"0041";
    tmp(49709) := x"0041";
    tmp(49710) := x"0041";
    tmp(49711) := x"0041";
    tmp(49712) := x"0061";
    tmp(49713) := x"0861";
    tmp(49714) := x"0862";
    tmp(49715) := x"0041";
    tmp(49716) := x"0041";
    tmp(49717) := x"0041";
    tmp(49718) := x"0021";
    tmp(49719) := x"0020";
    tmp(49720) := x"0020";
    tmp(49721) := x"0020";
    tmp(49722) := x"0020";
    tmp(49723) := x"0020";
    tmp(49724) := x"0000";
    tmp(49725) := x"0000";
    tmp(49726) := x"0000";
    tmp(49727) := x"0000";
    tmp(49728) := x"0000";
    tmp(49729) := x"0000";
    tmp(49730) := x"0000";
    tmp(49731) := x"0020";
    tmp(49732) := x"0020";
    tmp(49733) := x"0020";
    tmp(49734) := x"0020";
    tmp(49735) := x"0020";
    tmp(49736) := x"0020";
    tmp(49737) := x"0020";
    tmp(49738) := x"0020";
    tmp(49739) := x"0020";
    tmp(49740) := x"0020";
    tmp(49741) := x"0020";
    tmp(49742) := x"0021";
    tmp(49743) := x"0041";
    tmp(49744) := x"0041";
    tmp(49745) := x"0861";
    tmp(49746) := x"0862";
    tmp(49747) := x"0862";
    tmp(49748) := x"0882";
    tmp(49749) := x"08a3";
    tmp(49750) := x"08a3";
    tmp(49751) := x"08c4";
    tmp(49752) := x"08a3";
    tmp(49753) := x"08a3";
    tmp(49754) := x"0841";
    tmp(49755) := x"0820";
    tmp(49756) := x"1020";
    tmp(49757) := x"1020";
    tmp(49758) := x"1020";
    tmp(49759) := x"0840";
    tmp(49760) := x"0840";
    tmp(49761) := x"0820";
    tmp(49762) := x"0820";
    tmp(49763) := x"0820";
    tmp(49764) := x"0820";
    tmp(49765) := x"0820";
    tmp(49766) := x"0841";
    tmp(49767) := x"1061";
    tmp(49768) := x"1061";
    tmp(49769) := x"1041";
    tmp(49770) := x"1020";
    tmp(49771) := x"1020";
    tmp(49772) := x"1840";
    tmp(49773) := x"2061";
    tmp(49774) := x"1881";
    tmp(49775) := x"1880";
    tmp(49776) := x"2080";
    tmp(49777) := x"2081";
    tmp(49778) := x"28a1";
    tmp(49779) := x"28a1";
    tmp(49780) := x"2081";
    tmp(49781) := x"1861";
    tmp(49782) := x"1860";
    tmp(49783) := x"1060";
    tmp(49784) := x"1060";
    tmp(49785) := x"1060";
    tmp(49786) := x"1060";
    tmp(49787) := x"1060";
    tmp(49788) := x"1060";
    tmp(49789) := x"1060";
    tmp(49790) := x"0840";
    tmp(49791) := x"0840";
    tmp(49792) := x"0000";
    tmp(49793) := x"0000";
    tmp(49794) := x"0000";
    tmp(49795) := x"0000";
    tmp(49796) := x"0000";
    tmp(49797) := x"0000";
    tmp(49798) := x"0020";
    tmp(49799) := x"0000";
    tmp(49800) := x"0000";
    tmp(49801) := x"0000";
    tmp(49802) := x"0000";
    tmp(49803) := x"0000";
    tmp(49804) := x"0000";
    tmp(49805) := x"0000";
    tmp(49806) := x"0020";
    tmp(49807) := x"0020";
    tmp(49808) := x"0821";
    tmp(49809) := x"0020";
    tmp(49810) := x"0020";
    tmp(49811) := x"0020";
    tmp(49812) := x"0020";
    tmp(49813) := x"0000";
    tmp(49814) := x"0000";
    tmp(49815) := x"0000";
    tmp(49816) := x"0000";
    tmp(49817) := x"0000";
    tmp(49818) := x"0841";
    tmp(49819) := x"28a2";
    tmp(49820) := x"5944";
    tmp(49821) := x"50e3";
    tmp(49822) := x"4862";
    tmp(49823) := x"3021";
    tmp(49824) := x"5082";
    tmp(49825) := x"a229";
    tmp(49826) := x"6966";
    tmp(49827) := x"c32e";
    tmp(49828) := x"89a8";
    tmp(49829) := x"68e4";
    tmp(49830) := x"68e4";
    tmp(49831) := x"91c8";
    tmp(49832) := x"c2cd";
    tmp(49833) := x"60c4";
    tmp(49834) := x"3841";
    tmp(49835) := x"b1e8";
    tmp(49836) := x"99ea";
    tmp(49837) := x"a24b";
    tmp(49838) := x"91c8";
    tmp(49839) := x"68e4";
    tmp(49840) := x"4861";
    tmp(49841) := x"3821";
    tmp(49842) := x"9945";
    tmp(49843) := x"ca09";
    tmp(49844) := x"5882";
    tmp(49845) := x"5882";
    tmp(49846) := x"4821";
    tmp(49847) := x"3800";
    tmp(49848) := x"3800";
    tmp(49849) := x"4000";
    tmp(49850) := x"5800";
    tmp(49851) := x"5800";
    tmp(49852) := x"6000";
    tmp(49853) := x"7000";
    tmp(49854) := x"8820";
    tmp(49855) := x"a020";
    tmp(49856) := x"a020";
    tmp(49857) := x"b820";
    tmp(49858) := x"e020";
    tmp(49859) := x"d820";
    tmp(49860) := x"a800";
    tmp(49861) := x"d020";
    tmp(49862) := x"c820";
    tmp(49863) := x"c020";
    tmp(49864) := x"e020";
    tmp(49865) := x"c820";
    tmp(49866) := x"e840";
    tmp(49867) := x"f861";
    tmp(49868) := x"7061";
    tmp(49869) := x"1840";
    tmp(49870) := x"0840";
    tmp(49871) := x"0840";
    tmp(49872) := x"0840";
    tmp(49873) := x"0840";
    tmp(49874) := x"0840";
    tmp(49875) := x"0840";
    tmp(49876) := x"0840";
    tmp(49877) := x"0840";
    tmp(49878) := x"0840";
    tmp(49879) := x"0840";
    tmp(49880) := x"0840";
    tmp(49881) := x"0840";
    tmp(49882) := x"0840";
    tmp(49883) := x"0840";
    tmp(49884) := x"0840";
    tmp(49885) := x"0840";
    tmp(49886) := x"0840";
    tmp(49887) := x"0840";
    tmp(49888) := x"0840";
    tmp(49889) := x"0840";
    tmp(49890) := x"0840";
    tmp(49891) := x"0840";
    tmp(49892) := x"0840";
    tmp(49893) := x"0840";
    tmp(49894) := x"0840";
    tmp(49895) := x"0840";
    tmp(49896) := x"0840";
    tmp(49897) := x"0840";
    tmp(49898) := x"0840";
    tmp(49899) := x"0840";
    tmp(49900) := x"0840";
    tmp(49901) := x"0840";
    tmp(49902) := x"0840";
    tmp(49903) := x"0841";
    tmp(49904) := x"0840";
    tmp(49905) := x"0840";
    tmp(49906) := x"0840";
    tmp(49907) := x"0840";
    tmp(49908) := x"0840";
    tmp(49909) := x"0840";
    tmp(49910) := x"0840";
    tmp(49911) := x"0840";
    tmp(49912) := x"0840";
    tmp(49913) := x"0840";
    tmp(49914) := x"0840";
    tmp(49915) := x"0840";
    tmp(49916) := x"0840";
    tmp(49917) := x"0840";
    tmp(49918) := x"0840";
    tmp(49919) := x"0840";
    tmp(49920) := x"0000";
    tmp(49921) := x"08a0";
    tmp(49922) := x"08a0";
    tmp(49923) := x"08c0";
    tmp(49924) := x"08c0";
    tmp(49925) := x"08c0";
    tmp(49926) := x"08c0";
    tmp(49927) := x"08c0";
    tmp(49928) := x"08c0";
    tmp(49929) := x"08e1";
    tmp(49930) := x"08e1";
    tmp(49931) := x"08e1";
    tmp(49932) := x"08e1";
    tmp(49933) := x"10e1";
    tmp(49934) := x"10e1";
    tmp(49935) := x"1101";
    tmp(49936) := x"1101";
    tmp(49937) := x"1101";
    tmp(49938) := x"1101";
    tmp(49939) := x"08e1";
    tmp(49940) := x"08c2";
    tmp(49941) := x"0881";
    tmp(49942) := x"0061";
    tmp(49943) := x"0041";
    tmp(49944) := x"0041";
    tmp(49945) := x"0041";
    tmp(49946) := x"0041";
    tmp(49947) := x"0041";
    tmp(49948) := x"0841";
    tmp(49949) := x"0841";
    tmp(49950) := x"0841";
    tmp(49951) := x"0021";
    tmp(49952) := x"0020";
    tmp(49953) := x"0000";
    tmp(49954) := x"0000";
    tmp(49955) := x"0000";
    tmp(49956) := x"0000";
    tmp(49957) := x"0000";
    tmp(49958) := x"0000";
    tmp(49959) := x"0000";
    tmp(49960) := x"0000";
    tmp(49961) := x"0000";
    tmp(49962) := x"0000";
    tmp(49963) := x"0000";
    tmp(49964) := x"0000";
    tmp(49965) := x"0000";
    tmp(49966) := x"0000";
    tmp(49967) := x"0000";
    tmp(49968) := x"0800";
    tmp(49969) := x"0800";
    tmp(49970) := x"0800";
    tmp(49971) := x"0800";
    tmp(49972) := x"0800";
    tmp(49973) := x"0800";
    tmp(49974) := x"0800";
    tmp(49975) := x"0800";
    tmp(49976) := x"0800";
    tmp(49977) := x"0800";
    tmp(49978) := x"0000";
    tmp(49979) := x"0000";
    tmp(49980) := x"0800";
    tmp(49981) := x"0800";
    tmp(49982) := x"0820";
    tmp(49983) := x"0820";
    tmp(49984) := x"0820";
    tmp(49985) := x"0820";
    tmp(49986) := x"1041";
    tmp(49987) := x"1861";
    tmp(49988) := x"1061";
    tmp(49989) := x"0841";
    tmp(49990) := x"0841";
    tmp(49991) := x"1082";
    tmp(49992) := x"1062";
    tmp(49993) := x"0841";
    tmp(49994) := x"0821";
    tmp(49995) := x"0800";
    tmp(49996) := x"0800";
    tmp(49997) := x"1020";
    tmp(49998) := x"1820";
    tmp(49999) := x"1840";
    tmp(50000) := x"1040";
    tmp(50001) := x"0840";
    tmp(50002) := x"0820";
    tmp(50003) := x"0820";
    tmp(50004) := x"0840";
    tmp(50005) := x"0841";
    tmp(50006) := x"0841";
    tmp(50007) := x"0841";
    tmp(50008) := x"0841";
    tmp(50009) := x"0841";
    tmp(50010) := x"1020";
    tmp(50011) := x"1820";
    tmp(50012) := x"1020";
    tmp(50013) := x"1020";
    tmp(50014) := x"1020";
    tmp(50015) := x"1020";
    tmp(50016) := x"1040";
    tmp(50017) := x"1840";
    tmp(50018) := x"1860";
    tmp(50019) := x"2061";
    tmp(50020) := x"2061";
    tmp(50021) := x"2061";
    tmp(50022) := x"2041";
    tmp(50023) := x"2040";
    tmp(50024) := x"2040";
    tmp(50025) := x"2040";
    tmp(50026) := x"1840";
    tmp(50027) := x"1060";
    tmp(50028) := x"1040";
    tmp(50029) := x"1040";
    tmp(50030) := x"1840";
    tmp(50031) := x"1040";
    tmp(50032) := x"0000";
    tmp(50033) := x"0000";
    tmp(50034) := x"0000";
    tmp(50035) := x"0000";
    tmp(50036) := x"0000";
    tmp(50037) := x"0000";
    tmp(50038) := x"0000";
    tmp(50039) := x"0000";
    tmp(50040) := x"0000";
    tmp(50041) := x"0000";
    tmp(50042) := x"0000";
    tmp(50043) := x"0000";
    tmp(50044) := x"0000";
    tmp(50045) := x"0020";
    tmp(50046) := x"0821";
    tmp(50047) := x"0841";
    tmp(50048) := x"0021";
    tmp(50049) := x"0000";
    tmp(50050) := x"0000";
    tmp(50051) := x"0020";
    tmp(50052) := x"0820";
    tmp(50053) := x"0821";
    tmp(50054) := x"0820";
    tmp(50055) := x"0020";
    tmp(50056) := x"0820";
    tmp(50057) := x"0820";
    tmp(50058) := x"5186";
    tmp(50059) := x"2862";
    tmp(50060) := x"3082";
    tmp(50061) := x"9a08";
    tmp(50062) := x"ca8b";
    tmp(50063) := x"60c3";
    tmp(50064) := x"7145";
    tmp(50065) := x"dbd1";
    tmp(50066) := x"89e9";
    tmp(50067) := x"cb0e";
    tmp(50068) := x"50a3";
    tmp(50069) := x"eb6f";
    tmp(50070) := x"7926";
    tmp(50071) := x"91c8";
    tmp(50072) := x"baac";
    tmp(50073) := x"db4e";
    tmp(50074) := x"68a3";
    tmp(50075) := x"4041";
    tmp(50076) := x"70e4";
    tmp(50077) := x"aa4a";
    tmp(50078) := x"7104";
    tmp(50079) := x"4861";
    tmp(50080) := x"6082";
    tmp(50081) := x"4841";
    tmp(50082) := x"3000";
    tmp(50083) := x"5862";
    tmp(50084) := x"e28a";
    tmp(50085) := x"6062";
    tmp(50086) := x"3000";
    tmp(50087) := x"3800";
    tmp(50088) := x"4000";
    tmp(50089) := x"4800";
    tmp(50090) := x"5800";
    tmp(50091) := x"5800";
    tmp(50092) := x"6000";
    tmp(50093) := x"6800";
    tmp(50094) := x"8000";
    tmp(50095) := x"9000";
    tmp(50096) := x"9800";
    tmp(50097) := x"a800";
    tmp(50098) := x"d820";
    tmp(50099) := x"b000";
    tmp(50100) := x"a000";
    tmp(50101) := x"d820";
    tmp(50102) := x"c020";
    tmp(50103) := x"b820";
    tmp(50104) := x"e020";
    tmp(50105) := x"e040";
    tmp(50106) := x"f040";
    tmp(50107) := x"f861";
    tmp(50108) := x"6060";
    tmp(50109) := x"1040";
    tmp(50110) := x"0840";
    tmp(50111) := x"0840";
    tmp(50112) := x"0840";
    tmp(50113) := x"0840";
    tmp(50114) := x"0840";
    tmp(50115) := x"0840";
    tmp(50116) := x"0840";
    tmp(50117) := x"0840";
    tmp(50118) := x"0840";
    tmp(50119) := x"0840";
    tmp(50120) := x"0840";
    tmp(50121) := x"0840";
    tmp(50122) := x"0840";
    tmp(50123) := x"0840";
    tmp(50124) := x"0840";
    tmp(50125) := x"0840";
    tmp(50126) := x"0840";
    tmp(50127) := x"0840";
    tmp(50128) := x"0840";
    tmp(50129) := x"0840";
    tmp(50130) := x"0840";
    tmp(50131) := x"0840";
    tmp(50132) := x"0840";
    tmp(50133) := x"0840";
    tmp(50134) := x"0840";
    tmp(50135) := x"0840";
    tmp(50136) := x"0840";
    tmp(50137) := x"0840";
    tmp(50138) := x"0840";
    tmp(50139) := x"0840";
    tmp(50140) := x"0840";
    tmp(50141) := x"0840";
    tmp(50142) := x"0840";
    tmp(50143) := x"0840";
    tmp(50144) := x"0840";
    tmp(50145) := x"0840";
    tmp(50146) := x"0840";
    tmp(50147) := x"0840";
    tmp(50148) := x"0840";
    tmp(50149) := x"0840";
    tmp(50150) := x"0840";
    tmp(50151) := x"0840";
    tmp(50152) := x"0840";
    tmp(50153) := x"0840";
    tmp(50154) := x"0840";
    tmp(50155) := x"0840";
    tmp(50156) := x"0840";
    tmp(50157) := x"0840";
    tmp(50158) := x"0840";
    tmp(50159) := x"0840";
    tmp(50160) := x"0000";
    tmp(50161) := x"08c0";
    tmp(50162) := x"08a0";
    tmp(50163) := x"08c0";
    tmp(50164) := x"08a0";
    tmp(50165) := x"08a0";
    tmp(50166) := x"08a0";
    tmp(50167) := x"08c0";
    tmp(50168) := x"08c0";
    tmp(50169) := x"08c1";
    tmp(50170) := x"08e1";
    tmp(50171) := x"08e1";
    tmp(50172) := x"08e1";
    tmp(50173) := x"08e1";
    tmp(50174) := x"08e1";
    tmp(50175) := x"08c1";
    tmp(50176) := x"08c1";
    tmp(50177) := x"08a1";
    tmp(50178) := x"0881";
    tmp(50179) := x"0041";
    tmp(50180) := x"0021";
    tmp(50181) := x"0020";
    tmp(50182) := x"0021";
    tmp(50183) := x"0041";
    tmp(50184) := x"0821";
    tmp(50185) := x"0821";
    tmp(50186) := x"0821";
    tmp(50187) := x"0020";
    tmp(50188) := x"0000";
    tmp(50189) := x"0000";
    tmp(50190) := x"0000";
    tmp(50191) := x"0000";
    tmp(50192) := x"0000";
    tmp(50193) := x"0000";
    tmp(50194) := x"0000";
    tmp(50195) := x"0000";
    tmp(50196) := x"0800";
    tmp(50197) := x"0800";
    tmp(50198) := x"0800";
    tmp(50199) := x"0800";
    tmp(50200) := x"1000";
    tmp(50201) := x"1000";
    tmp(50202) := x"1000";
    tmp(50203) := x"1000";
    tmp(50204) := x"1800";
    tmp(50205) := x"1800";
    tmp(50206) := x"1800";
    tmp(50207) := x"1800";
    tmp(50208) := x"1800";
    tmp(50209) := x"1800";
    tmp(50210) := x"1800";
    tmp(50211) := x"1800";
    tmp(50212) := x"1800";
    tmp(50213) := x"1800";
    tmp(50214) := x"1800";
    tmp(50215) := x"2000";
    tmp(50216) := x"2000";
    tmp(50217) := x"2020";
    tmp(50218) := x"2020";
    tmp(50219) := x"2020";
    tmp(50220) := x"2020";
    tmp(50221) := x"2020";
    tmp(50222) := x"2020";
    tmp(50223) := x"1820";
    tmp(50224) := x"2020";
    tmp(50225) := x"2020";
    tmp(50226) := x"2020";
    tmp(50227) := x"2020";
    tmp(50228) := x"2020";
    tmp(50229) := x"2020";
    tmp(50230) := x"1820";
    tmp(50231) := x"1820";
    tmp(50232) := x"2041";
    tmp(50233) := x"2041";
    tmp(50234) := x"1820";
    tmp(50235) := x"1020";
    tmp(50236) := x"0800";
    tmp(50237) := x"0800";
    tmp(50238) := x"0800";
    tmp(50239) := x"1020";
    tmp(50240) := x"1020";
    tmp(50241) := x"1020";
    tmp(50242) := x"1020";
    tmp(50243) := x"0820";
    tmp(50244) := x"0820";
    tmp(50245) := x"0820";
    tmp(50246) := x"0841";
    tmp(50247) := x"0841";
    tmp(50248) := x"0841";
    tmp(50249) := x"0800";
    tmp(50250) := x"1020";
    tmp(50251) := x"1820";
    tmp(50252) := x"2020";
    tmp(50253) := x"1020";
    tmp(50254) := x"0800";
    tmp(50255) := x"0820";
    tmp(50256) := x"2040";
    tmp(50257) := x"3040";
    tmp(50258) := x"2820";
    tmp(50259) := x"2840";
    tmp(50260) := x"2841";
    tmp(50261) := x"2861";
    tmp(50262) := x"2041";
    tmp(50263) := x"2040";
    tmp(50264) := x"2820";
    tmp(50265) := x"3040";
    tmp(50266) := x"3040";
    tmp(50267) := x"2840";
    tmp(50268) := x"2840";
    tmp(50269) := x"2840";
    tmp(50270) := x"3040";
    tmp(50271) := x"2020";
    tmp(50272) := x"0000";
    tmp(50273) := x"0000";
    tmp(50274) := x"0000";
    tmp(50275) := x"0000";
    tmp(50276) := x"0000";
    tmp(50277) := x"0020";
    tmp(50278) := x"0020";
    tmp(50279) := x"0000";
    tmp(50280) := x"0000";
    tmp(50281) := x"0000";
    tmp(50282) := x"0000";
    tmp(50283) := x"0000";
    tmp(50284) := x"0000";
    tmp(50285) := x"0000";
    tmp(50286) := x"0000";
    tmp(50287) := x"0000";
    tmp(50288) := x"0020";
    tmp(50289) := x"0000";
    tmp(50290) := x"0000";
    tmp(50291) := x"0000";
    tmp(50292) := x"0020";
    tmp(50293) := x"0000";
    tmp(50294) := x"0821";
    tmp(50295) := x"0821";
    tmp(50296) := x"1041";
    tmp(50297) := x"2082";
    tmp(50298) := x"8249";
    tmp(50299) := x"48e4";
    tmp(50300) := x"40a2";
    tmp(50301) := x"9165";
    tmp(50302) := x"5062";
    tmp(50303) := x"4841";
    tmp(50304) := x"b26a";
    tmp(50305) := x"aa4a";
    tmp(50306) := x"bb0d";
    tmp(50307) := x"8987";
    tmp(50308) := x"60e4";
    tmp(50309) := x"ebd1";
    tmp(50310) := x"7105";
    tmp(50311) := x"89a7";
    tmp(50312) := x"7146";
    tmp(50313) := x"c2ac";
    tmp(50314) := x"68e4";
    tmp(50315) := x"78e4";
    tmp(50316) := x"4862";
    tmp(50317) := x"3841";
    tmp(50318) := x"5062";
    tmp(50319) := x"68a3";
    tmp(50320) := x"5882";
    tmp(50321) := x"4841";
    tmp(50322) := x"90c3";
    tmp(50323) := x"3000";
    tmp(50324) := x"5841";
    tmp(50325) := x"5841";
    tmp(50326) := x"2800";
    tmp(50327) := x"3800";
    tmp(50328) := x"4000";
    tmp(50329) := x"5000";
    tmp(50330) := x"5800";
    tmp(50331) := x"6000";
    tmp(50332) := x"6000";
    tmp(50333) := x"6800";
    tmp(50334) := x"8000";
    tmp(50335) := x"9000";
    tmp(50336) := x"9800";
    tmp(50337) := x"b020";
    tmp(50338) := x"d820";
    tmp(50339) := x"b000";
    tmp(50340) := x"a800";
    tmp(50341) := x"c820";
    tmp(50342) := x"c020";
    tmp(50343) := x"b000";
    tmp(50344) := x"c020";
    tmp(50345) := x"f841";
    tmp(50346) := x"e840";
    tmp(50347) := x"f861";
    tmp(50348) := x"5860";
    tmp(50349) := x"1040";
    tmp(50350) := x"0840";
    tmp(50351) := x"0840";
    tmp(50352) := x"0840";
    tmp(50353) := x"0840";
    tmp(50354) := x"0840";
    tmp(50355) := x"0840";
    tmp(50356) := x"0840";
    tmp(50357) := x"0840";
    tmp(50358) := x"0840";
    tmp(50359) := x"0840";
    tmp(50360) := x"0840";
    tmp(50361) := x"0840";
    tmp(50362) := x"0840";
    tmp(50363) := x"0840";
    tmp(50364) := x"0840";
    tmp(50365) := x"0840";
    tmp(50366) := x"0840";
    tmp(50367) := x"0840";
    tmp(50368) := x"0840";
    tmp(50369) := x"0840";
    tmp(50370) := x"0840";
    tmp(50371) := x"0840";
    tmp(50372) := x"0840";
    tmp(50373) := x"0840";
    tmp(50374) := x"0840";
    tmp(50375) := x"0840";
    tmp(50376) := x"0840";
    tmp(50377) := x"0840";
    tmp(50378) := x"0840";
    tmp(50379) := x"0840";
    tmp(50380) := x"0840";
    tmp(50381) := x"0840";
    tmp(50382) := x"0840";
    tmp(50383) := x"0840";
    tmp(50384) := x"0840";
    tmp(50385) := x"0840";
    tmp(50386) := x"0840";
    tmp(50387) := x"0840";
    tmp(50388) := x"0840";
    tmp(50389) := x"0840";
    tmp(50390) := x"0840";
    tmp(50391) := x"0840";
    tmp(50392) := x"0840";
    tmp(50393) := x"0840";
    tmp(50394) := x"0840";
    tmp(50395) := x"0840";
    tmp(50396) := x"0840";
    tmp(50397) := x"0840";
    tmp(50398) := x"0840";
    tmp(50399) := x"0840";
    tmp(50400) := x"0020";
    tmp(50401) := x"08c1";
    tmp(50402) := x"08c0";
    tmp(50403) := x"08c1";
    tmp(50404) := x"08c0";
    tmp(50405) := x"08a0";
    tmp(50406) := x"08a0";
    tmp(50407) := x"08a0";
    tmp(50408) := x"08c0";
    tmp(50409) := x"08c1";
    tmp(50410) := x"08c1";
    tmp(50411) := x"08c1";
    tmp(50412) := x"08a1";
    tmp(50413) := x"0881";
    tmp(50414) := x"0881";
    tmp(50415) := x"0061";
    tmp(50416) := x"0041";
    tmp(50417) := x"0020";
    tmp(50418) := x"0020";
    tmp(50419) := x"0020";
    tmp(50420) := x"0020";
    tmp(50421) := x"0821";
    tmp(50422) := x"0820";
    tmp(50423) := x"0820";
    tmp(50424) := x"0000";
    tmp(50425) := x"0000";
    tmp(50426) := x"0000";
    tmp(50427) := x"0000";
    tmp(50428) := x"0000";
    tmp(50429) := x"0000";
    tmp(50430) := x"0000";
    tmp(50431) := x"0000";
    tmp(50432) := x"0800";
    tmp(50433) := x"0800";
    tmp(50434) := x"0800";
    tmp(50435) := x"1000";
    tmp(50436) := x"1000";
    tmp(50437) := x"1800";
    tmp(50438) := x"1800";
    tmp(50439) := x"1800";
    tmp(50440) := x"1800";
    tmp(50441) := x"1800";
    tmp(50442) := x"1000";
    tmp(50443) := x"1000";
    tmp(50444) := x"1800";
    tmp(50445) := x"1800";
    tmp(50446) := x"1800";
    tmp(50447) := x"1800";
    tmp(50448) := x"1820";
    tmp(50449) := x"1820";
    tmp(50450) := x"1800";
    tmp(50451) := x"1800";
    tmp(50452) := x"1800";
    tmp(50453) := x"1800";
    tmp(50454) := x"2000";
    tmp(50455) := x"2020";
    tmp(50456) := x"2020";
    tmp(50457) := x"2820";
    tmp(50458) := x"2820";
    tmp(50459) := x"2840";
    tmp(50460) := x"2820";
    tmp(50461) := x"2820";
    tmp(50462) := x"2020";
    tmp(50463) := x"2000";
    tmp(50464) := x"1800";
    tmp(50465) := x"1800";
    tmp(50466) := x"1800";
    tmp(50467) := x"1820";
    tmp(50468) := x"2020";
    tmp(50469) := x"2020";
    tmp(50470) := x"2840";
    tmp(50471) := x"2840";
    tmp(50472) := x"3041";
    tmp(50473) := x"3041";
    tmp(50474) := x"3040";
    tmp(50475) := x"3041";
    tmp(50476) := x"2841";
    tmp(50477) := x"1821";
    tmp(50478) := x"1020";
    tmp(50479) := x"1020";
    tmp(50480) := x"0800";
    tmp(50481) := x"0800";
    tmp(50482) := x"1000";
    tmp(50483) := x"1000";
    tmp(50484) := x"0800";
    tmp(50485) := x"0800";
    tmp(50486) := x"0820";
    tmp(50487) := x"1020";
    tmp(50488) := x"1020";
    tmp(50489) := x"0800";
    tmp(50490) := x"0800";
    tmp(50491) := x"1000";
    tmp(50492) := x"1820";
    tmp(50493) := x"1000";
    tmp(50494) := x"0800";
    tmp(50495) := x"0820";
    tmp(50496) := x"1820";
    tmp(50497) := x"4020";
    tmp(50498) := x"4820";
    tmp(50499) := x"4820";
    tmp(50500) := x"4820";
    tmp(50501) := x"4020";
    tmp(50502) := x"4041";
    tmp(50503) := x"3020";
    tmp(50504) := x"2820";
    tmp(50505) := x"3020";
    tmp(50506) := x"4040";
    tmp(50507) := x"4820";
    tmp(50508) := x"3820";
    tmp(50509) := x"3820";
    tmp(50510) := x"3820";
    tmp(50511) := x"2020";
    tmp(50512) := x"0000";
    tmp(50513) := x"0000";
    tmp(50514) := x"0000";
    tmp(50515) := x"0000";
    tmp(50516) := x"0000";
    tmp(50517) := x"0000";
    tmp(50518) := x"0020";
    tmp(50519) := x"0000";
    tmp(50520) := x"0000";
    tmp(50521) := x"0000";
    tmp(50522) := x"0000";
    tmp(50523) := x"0000";
    tmp(50524) := x"0000";
    tmp(50525) := x"0000";
    tmp(50526) := x"0000";
    tmp(50527) := x"0000";
    tmp(50528) := x"0020";
    tmp(50529) := x"0000";
    tmp(50530) := x"0000";
    tmp(50531) := x"0020";
    tmp(50532) := x"0020";
    tmp(50533) := x"0000";
    tmp(50534) := x"0820";
    tmp(50535) := x"1062";
    tmp(50536) := x"0821";
    tmp(50537) := x"38e4";
    tmp(50538) := x"ab0d";
    tmp(50539) := x"58e4";
    tmp(50540) := x"58c3";
    tmp(50541) := x"5841";
    tmp(50542) := x"4020";
    tmp(50543) := x"6082";
    tmp(50544) := x"d34f";
    tmp(50545) := x"91e9";
    tmp(50546) := x"aa4a";
    tmp(50547) := x"58a3";
    tmp(50548) := x"c28a";
    tmp(50549) := x"d2ed";
    tmp(50550) := x"4882";
    tmp(50551) := x"b26a";
    tmp(50552) := x"68e4";
    tmp(50553) := x"8966";
    tmp(50554) := x"8126";
    tmp(50555) := x"58c4";
    tmp(50556) := x"cacc";
    tmp(50557) := x"8146";
    tmp(50558) := x"5082";
    tmp(50559) := x"4041";
    tmp(50560) := x"3841";
    tmp(50561) := x"5882";
    tmp(50562) := x"60a3";
    tmp(50563) := x"3820";
    tmp(50564) := x"2800";
    tmp(50565) := x"3820";
    tmp(50566) := x"3000";
    tmp(50567) := x"3800";
    tmp(50568) := x"4800";
    tmp(50569) := x"6820";
    tmp(50570) := x"6000";
    tmp(50571) := x"6000";
    tmp(50572) := x"5800";
    tmp(50573) := x"6800";
    tmp(50574) := x"8820";
    tmp(50575) := x"9000";
    tmp(50576) := x"a000";
    tmp(50577) := x"b000";
    tmp(50578) := x"c820";
    tmp(50579) := x"a000";
    tmp(50580) := x"a000";
    tmp(50581) := x"b820";
    tmp(50582) := x"b800";
    tmp(50583) := x"c020";
    tmp(50584) := x"b820";
    tmp(50585) := x"f040";
    tmp(50586) := x"e840";
    tmp(50587) := x"f861";
    tmp(50588) := x"6060";
    tmp(50589) := x"1040";
    tmp(50590) := x"0840";
    tmp(50591) := x"0840";
    tmp(50592) := x"0840";
    tmp(50593) := x"0840";
    tmp(50594) := x"0840";
    tmp(50595) := x"0840";
    tmp(50596) := x"0840";
    tmp(50597) := x"0840";
    tmp(50598) := x"0840";
    tmp(50599) := x"0840";
    tmp(50600) := x"0840";
    tmp(50601) := x"0840";
    tmp(50602) := x"0840";
    tmp(50603) := x"0840";
    tmp(50604) := x"0840";
    tmp(50605) := x"0840";
    tmp(50606) := x"0840";
    tmp(50607) := x"0840";
    tmp(50608) := x"0840";
    tmp(50609) := x"0840";
    tmp(50610) := x"0840";
    tmp(50611) := x"0840";
    tmp(50612) := x"0840";
    tmp(50613) := x"0840";
    tmp(50614) := x"0840";
    tmp(50615) := x"0840";
    tmp(50616) := x"0840";
    tmp(50617) := x"0840";
    tmp(50618) := x"0840";
    tmp(50619) := x"0840";
    tmp(50620) := x"0840";
    tmp(50621) := x"0840";
    tmp(50622) := x"0840";
    tmp(50623) := x"0840";
    tmp(50624) := x"0840";
    tmp(50625) := x"0840";
    tmp(50626) := x"0840";
    tmp(50627) := x"0840";
    tmp(50628) := x"0840";
    tmp(50629) := x"0840";
    tmp(50630) := x"0840";
    tmp(50631) := x"0840";
    tmp(50632) := x"0840";
    tmp(50633) := x"0840";
    tmp(50634) := x"0840";
    tmp(50635) := x"0840";
    tmp(50636) := x"0840";
    tmp(50637) := x"0840";
    tmp(50638) := x"0840";
    tmp(50639) := x"0840";
    tmp(50640) := x"0020";
    tmp(50641) := x"08c1";
    tmp(50642) := x"08c1";
    tmp(50643) := x"08c1";
    tmp(50644) := x"08c1";
    tmp(50645) := x"08c0";
    tmp(50646) := x"08a0";
    tmp(50647) := x"08a0";
    tmp(50648) := x"08a1";
    tmp(50649) := x"08a1";
    tmp(50650) := x"0860";
    tmp(50651) := x"0040";
    tmp(50652) := x"0020";
    tmp(50653) := x"0020";
    tmp(50654) := x"0020";
    tmp(50655) := x"0020";
    tmp(50656) := x"0000";
    tmp(50657) := x"0000";
    tmp(50658) := x"0820";
    tmp(50659) := x"0820";
    tmp(50660) := x"0800";
    tmp(50661) := x"0800";
    tmp(50662) := x"0000";
    tmp(50663) := x"0000";
    tmp(50664) := x"0000";
    tmp(50665) := x"0000";
    tmp(50666) := x"0000";
    tmp(50667) := x"0000";
    tmp(50668) := x"0800";
    tmp(50669) := x"0800";
    tmp(50670) := x"0800";
    tmp(50671) := x"0800";
    tmp(50672) := x"1000";
    tmp(50673) := x"1000";
    tmp(50674) := x"1000";
    tmp(50675) := x"1000";
    tmp(50676) := x"1000";
    tmp(50677) := x"1800";
    tmp(50678) := x"1800";
    tmp(50679) := x"1800";
    tmp(50680) := x"1820";
    tmp(50681) := x"1820";
    tmp(50682) := x"1000";
    tmp(50683) := x"1000";
    tmp(50684) := x"1000";
    tmp(50685) := x"1000";
    tmp(50686) := x"1000";
    tmp(50687) := x"1000";
    tmp(50688) := x"1020";
    tmp(50689) := x"1020";
    tmp(50690) := x"1000";
    tmp(50691) := x"1000";
    tmp(50692) := x"1000";
    tmp(50693) := x"1000";
    tmp(50694) := x"1020";
    tmp(50695) := x"1820";
    tmp(50696) := x"1820";
    tmp(50697) := x"1820";
    tmp(50698) := x"1820";
    tmp(50699) := x"1820";
    tmp(50700) := x"1020";
    tmp(50701) := x"1000";
    tmp(50702) := x"1000";
    tmp(50703) := x"1000";
    tmp(50704) := x"1000";
    tmp(50705) := x"1000";
    tmp(50706) := x"1020";
    tmp(50707) := x"1020";
    tmp(50708) := x"1020";
    tmp(50709) := x"1020";
    tmp(50710) := x"1020";
    tmp(50711) := x"1020";
    tmp(50712) := x"1820";
    tmp(50713) := x"1840";
    tmp(50714) := x"2020";
    tmp(50715) := x"2040";
    tmp(50716) := x"2041";
    tmp(50717) := x"2041";
    tmp(50718) := x"1820";
    tmp(50719) := x"1820";
    tmp(50720) := x"2020";
    tmp(50721) := x"1800";
    tmp(50722) := x"1800";
    tmp(50723) := x"1800";
    tmp(50724) := x"1000";
    tmp(50725) := x"1000";
    tmp(50726) := x"1800";
    tmp(50727) := x"1820";
    tmp(50728) := x"1800";
    tmp(50729) := x"1800";
    tmp(50730) := x"1000";
    tmp(50731) := x"1000";
    tmp(50732) := x"2020";
    tmp(50733) := x"1820";
    tmp(50734) := x"0800";
    tmp(50735) := x"1020";
    tmp(50736) := x"2820";
    tmp(50737) := x"3820";
    tmp(50738) := x"4020";
    tmp(50739) := x"5020";
    tmp(50740) := x"5020";
    tmp(50741) := x"4820";
    tmp(50742) := x"4020";
    tmp(50743) := x"4020";
    tmp(50744) := x"4020";
    tmp(50745) := x"3820";
    tmp(50746) := x"3820";
    tmp(50747) := x"3820";
    tmp(50748) := x"3020";
    tmp(50749) := x"3020";
    tmp(50750) := x"3020";
    tmp(50751) := x"1800";
    tmp(50752) := x"0000";
    tmp(50753) := x"0000";
    tmp(50754) := x"0000";
    tmp(50755) := x"0000";
    tmp(50756) := x"0000";
    tmp(50757) := x"0000";
    tmp(50758) := x"0000";
    tmp(50759) := x"0000";
    tmp(50760) := x"0000";
    tmp(50761) := x"0000";
    tmp(50762) := x"0000";
    tmp(50763) := x"0000";
    tmp(50764) := x"0000";
    tmp(50765) := x"0000";
    tmp(50766) := x"0000";
    tmp(50767) := x"0000";
    tmp(50768) := x"0000";
    tmp(50769) := x"0000";
    tmp(50770) := x"0000";
    tmp(50771) := x"0020";
    tmp(50772) := x"0020";
    tmp(50773) := x"0000";
    tmp(50774) := x"0000";
    tmp(50775) := x"0841";
    tmp(50776) := x"1021";
    tmp(50777) := x"8a6a";
    tmp(50778) := x"9a8b";
    tmp(50779) := x"50c3";
    tmp(50780) := x"8925";
    tmp(50781) := x"6882";
    tmp(50782) := x"5861";
    tmp(50783) := x"8125";
    tmp(50784) := x"b26a";
    tmp(50785) := x"8187";
    tmp(50786) := x"aa09";
    tmp(50787) := x"4862";
    tmp(50788) := x"cb0d";
    tmp(50789) := x"e34f";
    tmp(50790) := x"4062";
    tmp(50791) := x"eb90";
    tmp(50792) := x"68c3";
    tmp(50793) := x"7125";
    tmp(50794) := x"91a8";
    tmp(50795) := x"6925";
    tmp(50796) := x"b28c";
    tmp(50797) := x"6925";
    tmp(50798) := x"91c8";
    tmp(50799) := x"9186";
    tmp(50800) := x"4041";
    tmp(50801) := x"4042";
    tmp(50802) := x"70c3";
    tmp(50803) := x"68a2";
    tmp(50804) := x"3020";
    tmp(50805) := x"3020";
    tmp(50806) := x"3000";
    tmp(50807) := x"4000";
    tmp(50808) := x"4800";
    tmp(50809) := x"6820";
    tmp(50810) := x"7000";
    tmp(50811) := x"6800";
    tmp(50812) := x"5800";
    tmp(50813) := x"7000";
    tmp(50814) := x"8800";
    tmp(50815) := x"9000";
    tmp(50816) := x"a800";
    tmp(50817) := x"a800";
    tmp(50818) := x"c020";
    tmp(50819) := x"a000";
    tmp(50820) := x"9800";
    tmp(50821) := x"b020";
    tmp(50822) := x"b000";
    tmp(50823) := x"c820";
    tmp(50824) := x"c020";
    tmp(50825) := x"e840";
    tmp(50826) := x"e840";
    tmp(50827) := x"f881";
    tmp(50828) := x"5860";
    tmp(50829) := x"1040";
    tmp(50830) := x"0840";
    tmp(50831) := x"0840";
    tmp(50832) := x"0840";
    tmp(50833) := x"0840";
    tmp(50834) := x"0840";
    tmp(50835) := x"0840";
    tmp(50836) := x"0840";
    tmp(50837) := x"0840";
    tmp(50838) := x"0840";
    tmp(50839) := x"0840";
    tmp(50840) := x"0840";
    tmp(50841) := x"0840";
    tmp(50842) := x"0840";
    tmp(50843) := x"0840";
    tmp(50844) := x"0840";
    tmp(50845) := x"0840";
    tmp(50846) := x"0840";
    tmp(50847) := x"0840";
    tmp(50848) := x"0840";
    tmp(50849) := x"0840";
    tmp(50850) := x"0840";
    tmp(50851) := x"0840";
    tmp(50852) := x"0840";
    tmp(50853) := x"0840";
    tmp(50854) := x"0840";
    tmp(50855) := x"0840";
    tmp(50856) := x"0840";
    tmp(50857) := x"0840";
    tmp(50858) := x"0840";
    tmp(50859) := x"0841";
    tmp(50860) := x"0840";
    tmp(50861) := x"0840";
    tmp(50862) := x"0840";
    tmp(50863) := x"0840";
    tmp(50864) := x"0840";
    tmp(50865) := x"0840";
    tmp(50866) := x"0840";
    tmp(50867) := x"0840";
    tmp(50868) := x"0840";
    tmp(50869) := x"0840";
    tmp(50870) := x"0840";
    tmp(50871) := x"0840";
    tmp(50872) := x"0840";
    tmp(50873) := x"0840";
    tmp(50874) := x"0840";
    tmp(50875) := x"0840";
    tmp(50876) := x"0840";
    tmp(50877) := x"0840";
    tmp(50878) := x"0840";
    tmp(50879) := x"0840";
    tmp(50880) := x"0020";
    tmp(50881) := x"08e1";
    tmp(50882) := x"08e1";
    tmp(50883) := x"08e1";
    tmp(50884) := x"08e1";
    tmp(50885) := x"08c1";
    tmp(50886) := x"08a1";
    tmp(50887) := x"0860";
    tmp(50888) := x"0040";
    tmp(50889) := x"0020";
    tmp(50890) := x"0020";
    tmp(50891) := x"0020";
    tmp(50892) := x"0000";
    tmp(50893) := x"0000";
    tmp(50894) := x"0000";
    tmp(50895) := x"0020";
    tmp(50896) := x"0820";
    tmp(50897) := x"0820";
    tmp(50898) := x"0800";
    tmp(50899) := x"0800";
    tmp(50900) := x"0000";
    tmp(50901) := x"0000";
    tmp(50902) := x"0000";
    tmp(50903) := x"0000";
    tmp(50904) := x"0000";
    tmp(50905) := x"0800";
    tmp(50906) := x"0800";
    tmp(50907) := x"0800";
    tmp(50908) := x"1000";
    tmp(50909) := x"1020";
    tmp(50910) := x"0800";
    tmp(50911) := x"0800";
    tmp(50912) := x"1000";
    tmp(50913) := x"1000";
    tmp(50914) := x"1000";
    tmp(50915) := x"1000";
    tmp(50916) := x"1000";
    tmp(50917) := x"1000";
    tmp(50918) := x"1000";
    tmp(50919) := x"1000";
    tmp(50920) := x"1020";
    tmp(50921) := x"1000";
    tmp(50922) := x"1000";
    tmp(50923) := x"1000";
    tmp(50924) := x"1000";
    tmp(50925) := x"1000";
    tmp(50926) := x"1000";
    tmp(50927) := x"1000";
    tmp(50928) := x"1000";
    tmp(50929) := x"1000";
    tmp(50930) := x"0800";
    tmp(50931) := x"1000";
    tmp(50932) := x"1000";
    tmp(50933) := x"1000";
    tmp(50934) := x"1020";
    tmp(50935) := x"1020";
    tmp(50936) := x"1020";
    tmp(50937) := x"1020";
    tmp(50938) := x"1020";
    tmp(50939) := x"1020";
    tmp(50940) := x"1000";
    tmp(50941) := x"1000";
    tmp(50942) := x"1000";
    tmp(50943) := x"0800";
    tmp(50944) := x"0800";
    tmp(50945) := x"0800";
    tmp(50946) := x"0820";
    tmp(50947) := x"0820";
    tmp(50948) := x"0820";
    tmp(50949) := x"0820";
    tmp(50950) := x"0820";
    tmp(50951) := x"0820";
    tmp(50952) := x"0820";
    tmp(50953) := x"0820";
    tmp(50954) := x"1020";
    tmp(50955) := x"1020";
    tmp(50956) := x"1020";
    tmp(50957) := x"1820";
    tmp(50958) := x"2020";
    tmp(50959) := x"2820";
    tmp(50960) := x"3020";
    tmp(50961) := x"3820";
    tmp(50962) := x"4020";
    tmp(50963) := x"4020";
    tmp(50964) := x"4020";
    tmp(50965) := x"4020";
    tmp(50966) := x"4040";
    tmp(50967) := x"4840";
    tmp(50968) := x"4841";
    tmp(50969) := x"4841";
    tmp(50970) := x"3841";
    tmp(50971) := x"3841";
    tmp(50972) := x"3841";
    tmp(50973) := x"3841";
    tmp(50974) := x"2020";
    tmp(50975) := x"2820";
    tmp(50976) := x"3820";
    tmp(50977) := x"3000";
    tmp(50978) := x"3820";
    tmp(50979) := x"4820";
    tmp(50980) := x"4820";
    tmp(50981) := x"4020";
    tmp(50982) := x"3820";
    tmp(50983) := x"3820";
    tmp(50984) := x"3820";
    tmp(50985) := x"3820";
    tmp(50986) := x"2820";
    tmp(50987) := x"2020";
    tmp(50988) := x"2000";
    tmp(50989) := x"2000";
    tmp(50990) := x"2000";
    tmp(50991) := x"1000";
    tmp(50992) := x"0000";
    tmp(50993) := x"0000";
    tmp(50994) := x"0000";
    tmp(50995) := x"0000";
    tmp(50996) := x"0000";
    tmp(50997) := x"0000";
    tmp(50998) := x"0000";
    tmp(50999) := x"0000";
    tmp(51000) := x"0000";
    tmp(51001) := x"0000";
    tmp(51002) := x"0000";
    tmp(51003) := x"0000";
    tmp(51004) := x"0000";
    tmp(51005) := x"0000";
    tmp(51006) := x"0000";
    tmp(51007) := x"0000";
    tmp(51008) := x"0000";
    tmp(51009) := x"0000";
    tmp(51010) := x"0000";
    tmp(51011) := x"0000";
    tmp(51012) := x"0020";
    tmp(51013) := x"0000";
    tmp(51014) := x"0000";
    tmp(51015) := x"0821";
    tmp(51016) := x"69c7";
    tmp(51017) := x"cbb1";
    tmp(51018) := x"6145";
    tmp(51019) := x"5904";
    tmp(51020) := x"e32e";
    tmp(51021) := x"c26b";
    tmp(51022) := x"9187";
    tmp(51023) := x"ba8b";
    tmp(51024) := x"6946";
    tmp(51025) := x"aa6a";
    tmp(51026) := x"60e4";
    tmp(51027) := x"8987";
    tmp(51028) := x"b26b";
    tmp(51029) := x"7926";
    tmp(51030) := x"5082";
    tmp(51031) := x"eb6e";
    tmp(51032) := x"68c4";
    tmp(51033) := x"7125";
    tmp(51034) := x"9209";
    tmp(51035) := x"58e4";
    tmp(51036) := x"8187";
    tmp(51037) := x"89c8";
    tmp(51038) := x"9a6c";
    tmp(51039) := x"924c";
    tmp(51040) := x"89e9";
    tmp(51041) := x"81a7";
    tmp(51042) := x"ba6a";
    tmp(51043) := x"daab";
    tmp(51044) := x"9145";
    tmp(51045) := x"3000";
    tmp(51046) := x"3000";
    tmp(51047) := x"4800";
    tmp(51048) := x"5000";
    tmp(51049) := x"6000";
    tmp(51050) := x"7800";
    tmp(51051) := x"7800";
    tmp(51052) := x"6800";
    tmp(51053) := x"7800";
    tmp(51054) := x"8800";
    tmp(51055) := x"9000";
    tmp(51056) := x"9800";
    tmp(51057) := x"a000";
    tmp(51058) := x"b020";
    tmp(51059) := x"9800";
    tmp(51060) := x"9000";
    tmp(51061) := x"c020";
    tmp(51062) := x"b820";
    tmp(51063) := x"d020";
    tmp(51064) := x"c020";
    tmp(51065) := x"d820";
    tmp(51066) := x"f040";
    tmp(51067) := x"f881";
    tmp(51068) := x"5860";
    tmp(51069) := x"1020";
    tmp(51070) := x"0840";
    tmp(51071) := x"0840";
    tmp(51072) := x"0840";
    tmp(51073) := x"0840";
    tmp(51074) := x"0840";
    tmp(51075) := x"0840";
    tmp(51076) := x"0840";
    tmp(51077) := x"0840";
    tmp(51078) := x"0840";
    tmp(51079) := x"0840";
    tmp(51080) := x"0840";
    tmp(51081) := x"0840";
    tmp(51082) := x"0840";
    tmp(51083) := x"0840";
    tmp(51084) := x"0840";
    tmp(51085) := x"0840";
    tmp(51086) := x"0840";
    tmp(51087) := x"0840";
    tmp(51088) := x"0840";
    tmp(51089) := x"0840";
    tmp(51090) := x"0840";
    tmp(51091) := x"0840";
    tmp(51092) := x"0840";
    tmp(51093) := x"0840";
    tmp(51094) := x"0840";
    tmp(51095) := x"0840";
    tmp(51096) := x"0840";
    tmp(51097) := x"0840";
    tmp(51098) := x"0840";
    tmp(51099) := x"0840";
    tmp(51100) := x"0840";
    tmp(51101) := x"0840";
    tmp(51102) := x"0840";
    tmp(51103) := x"0840";
    tmp(51104) := x"0840";
    tmp(51105) := x"0840";
    tmp(51106) := x"0840";
    tmp(51107) := x"0840";
    tmp(51108) := x"0840";
    tmp(51109) := x"0840";
    tmp(51110) := x"0840";
    tmp(51111) := x"0840";
    tmp(51112) := x"0840";
    tmp(51113) := x"0840";
    tmp(51114) := x"0840";
    tmp(51115) := x"0840";
    tmp(51116) := x"0840";
    tmp(51117) := x"0840";
    tmp(51118) := x"0840";
    tmp(51119) := x"0840";
    tmp(51120) := x"0020";
    tmp(51121) := x"08e1";
    tmp(51122) := x"10e1";
    tmp(51123) := x"08e1";
    tmp(51124) := x"08a1";
    tmp(51125) := x"0860";
    tmp(51126) := x"0020";
    tmp(51127) := x"0020";
    tmp(51128) := x"0000";
    tmp(51129) := x"0000";
    tmp(51130) := x"0000";
    tmp(51131) := x"0000";
    tmp(51132) := x"0000";
    tmp(51133) := x"0000";
    tmp(51134) := x"0820";
    tmp(51135) := x"0820";
    tmp(51136) := x"0820";
    tmp(51137) := x"0000";
    tmp(51138) := x"0000";
    tmp(51139) := x"0000";
    tmp(51140) := x"0000";
    tmp(51141) := x"0000";
    tmp(51142) := x"0800";
    tmp(51143) := x"0800";
    tmp(51144) := x"0800";
    tmp(51145) := x"0800";
    tmp(51146) := x"1000";
    tmp(51147) := x"1000";
    tmp(51148) := x"1000";
    tmp(51149) := x"1020";
    tmp(51150) := x"0800";
    tmp(51151) := x"0800";
    tmp(51152) := x"0800";
    tmp(51153) := x"0800";
    tmp(51154) := x"0800";
    tmp(51155) := x"0800";
    tmp(51156) := x"1000";
    tmp(51157) := x"1000";
    tmp(51158) := x"1000";
    tmp(51159) := x"1000";
    tmp(51160) := x"1000";
    tmp(51161) := x"1000";
    tmp(51162) := x"1000";
    tmp(51163) := x"0800";
    tmp(51164) := x"1000";
    tmp(51165) := x"1000";
    tmp(51166) := x"1000";
    tmp(51167) := x"1000";
    tmp(51168) := x"1000";
    tmp(51169) := x"1000";
    tmp(51170) := x"0800";
    tmp(51171) := x"0800";
    tmp(51172) := x"0800";
    tmp(51173) := x"0800";
    tmp(51174) := x"1000";
    tmp(51175) := x"1000";
    tmp(51176) := x"1000";
    tmp(51177) := x"1000";
    tmp(51178) := x"1020";
    tmp(51179) := x"1020";
    tmp(51180) := x"0800";
    tmp(51181) := x"1000";
    tmp(51182) := x"0800";
    tmp(51183) := x"0800";
    tmp(51184) := x"0800";
    tmp(51185) := x"0800";
    tmp(51186) := x"0820";
    tmp(51187) := x"0820";
    tmp(51188) := x"0820";
    tmp(51189) := x"0820";
    tmp(51190) := x"0820";
    tmp(51191) := x"0820";
    tmp(51192) := x"0800";
    tmp(51193) := x"0800";
    tmp(51194) := x"0820";
    tmp(51195) := x"0800";
    tmp(51196) := x"0800";
    tmp(51197) := x"1020";
    tmp(51198) := x"2020";
    tmp(51199) := x"3020";
    tmp(51200) := x"3820";
    tmp(51201) := x"4020";
    tmp(51202) := x"4820";
    tmp(51203) := x"4020";
    tmp(51204) := x"4020";
    tmp(51205) := x"4020";
    tmp(51206) := x"4820";
    tmp(51207) := x"4840";
    tmp(51208) := x"5841";
    tmp(51209) := x"6061";
    tmp(51210) := x"6081";
    tmp(51211) := x"6081";
    tmp(51212) := x"5041";
    tmp(51213) := x"4020";
    tmp(51214) := x"4020";
    tmp(51215) := x"4020";
    tmp(51216) := x"3820";
    tmp(51217) := x"3000";
    tmp(51218) := x"3000";
    tmp(51219) := x"3820";
    tmp(51220) := x"4020";
    tmp(51221) := x"4020";
    tmp(51222) := x"3820";
    tmp(51223) := x"3020";
    tmp(51224) := x"3020";
    tmp(51225) := x"3020";
    tmp(51226) := x"2820";
    tmp(51227) := x"2020";
    tmp(51228) := x"1800";
    tmp(51229) := x"1800";
    tmp(51230) := x"1800";
    tmp(51231) := x"0800";
    tmp(51232) := x"0000";
    tmp(51233) := x"0000";
    tmp(51234) := x"0000";
    tmp(51235) := x"0000";
    tmp(51236) := x"0000";
    tmp(51237) := x"0000";
    tmp(51238) := x"0000";
    tmp(51239) := x"0000";
    tmp(51240) := x"0000";
    tmp(51241) := x"0000";
    tmp(51242) := x"0000";
    tmp(51243) := x"0000";
    tmp(51244) := x"0000";
    tmp(51245) := x"0000";
    tmp(51246) := x"0000";
    tmp(51247) := x"0000";
    tmp(51248) := x"0000";
    tmp(51249) := x"0000";
    tmp(51250) := x"0000";
    tmp(51251) := x"0000";
    tmp(51252) := x"0020";
    tmp(51253) := x"0000";
    tmp(51254) := x"0000";
    tmp(51255) := x"38c3";
    tmp(51256) := x"dbf1";
    tmp(51257) := x"8a0a";
    tmp(51258) := x"50e4";
    tmp(51259) := x"aa49";
    tmp(51260) := x"e390";
    tmp(51261) := x"9209";
    tmp(51262) := x"9a2a";
    tmp(51263) := x"cb4f";
    tmp(51264) := x"7987";
    tmp(51265) := x"b26a";
    tmp(51266) := x"50a3";
    tmp(51267) := x"cacc";
    tmp(51268) := x"7946";
    tmp(51269) := x"8946";
    tmp(51270) := x"8125";
    tmp(51271) := x"91e8";
    tmp(51272) := x"4882";
    tmp(51273) := x"91e8";
    tmp(51274) := x"926b";
    tmp(51275) := x"79c8";
    tmp(51276) := x"81e8";
    tmp(51277) := x"926b";
    tmp(51278) := x"92cd";
    tmp(51279) := x"9b30";
    tmp(51280) := x"92ee";
    tmp(51281) := x"69c8";
    tmp(51282) := x"7166";
    tmp(51283) := x"c28a";
    tmp(51284) := x"fbaf";
    tmp(51285) := x"5861";
    tmp(51286) := x"3000";
    tmp(51287) := x"4000";
    tmp(51288) := x"5000";
    tmp(51289) := x"6000";
    tmp(51290) := x"7800";
    tmp(51291) := x"7800";
    tmp(51292) := x"6800";
    tmp(51293) := x"6800";
    tmp(51294) := x"8000";
    tmp(51295) := x"9000";
    tmp(51296) := x"9000";
    tmp(51297) := x"a800";
    tmp(51298) := x"a800";
    tmp(51299) := x"9800";
    tmp(51300) := x"9800";
    tmp(51301) := x"c820";
    tmp(51302) := x"c020";
    tmp(51303) := x"c820";
    tmp(51304) := x"b820";
    tmp(51305) := x"d820";
    tmp(51306) := x"f061";
    tmp(51307) := x"f8a1";
    tmp(51308) := x"5840";
    tmp(51309) := x"1020";
    tmp(51310) := x"0840";
    tmp(51311) := x"0840";
    tmp(51312) := x"0840";
    tmp(51313) := x"0840";
    tmp(51314) := x"0840";
    tmp(51315) := x"0840";
    tmp(51316) := x"0840";
    tmp(51317) := x"0840";
    tmp(51318) := x"0840";
    tmp(51319) := x"0840";
    tmp(51320) := x"0840";
    tmp(51321) := x"0840";
    tmp(51322) := x"0840";
    tmp(51323) := x"0840";
    tmp(51324) := x"0840";
    tmp(51325) := x"0840";
    tmp(51326) := x"0840";
    tmp(51327) := x"0840";
    tmp(51328) := x"0840";
    tmp(51329) := x"0840";
    tmp(51330) := x"0840";
    tmp(51331) := x"0840";
    tmp(51332) := x"0840";
    tmp(51333) := x"0840";
    tmp(51334) := x"0840";
    tmp(51335) := x"0840";
    tmp(51336) := x"0840";
    tmp(51337) := x"0840";
    tmp(51338) := x"0840";
    tmp(51339) := x"0840";
    tmp(51340) := x"0840";
    tmp(51341) := x"0840";
    tmp(51342) := x"0840";
    tmp(51343) := x"0840";
    tmp(51344) := x"0840";
    tmp(51345) := x"0840";
    tmp(51346) := x"0840";
    tmp(51347) := x"0840";
    tmp(51348) := x"0840";
    tmp(51349) := x"0840";
    tmp(51350) := x"0840";
    tmp(51351) := x"0840";
    tmp(51352) := x"0840";
    tmp(51353) := x"0840";
    tmp(51354) := x"0840";
    tmp(51355) := x"0840";
    tmp(51356) := x"0840";
    tmp(51357) := x"0840";
    tmp(51358) := x"0840";
    tmp(51359) := x"0840";
    tmp(51360) := x"0020";
    tmp(51361) := x"10e1";
    tmp(51362) := x"08a1";
    tmp(51363) := x"0860";
    tmp(51364) := x"0020";
    tmp(51365) := x"0000";
    tmp(51366) := x"0000";
    tmp(51367) := x"0000";
    tmp(51368) := x"0000";
    tmp(51369) := x"0000";
    tmp(51370) := x"0000";
    tmp(51371) := x"0000";
    tmp(51372) := x"0820";
    tmp(51373) := x"0820";
    tmp(51374) := x"0820";
    tmp(51375) := x"0000";
    tmp(51376) := x"0000";
    tmp(51377) := x"0000";
    tmp(51378) := x"0000";
    tmp(51379) := x"0000";
    tmp(51380) := x"0000";
    tmp(51381) := x"0800";
    tmp(51382) := x"0800";
    tmp(51383) := x"0800";
    tmp(51384) := x"0800";
    tmp(51385) := x"0800";
    tmp(51386) := x"0800";
    tmp(51387) := x"1000";
    tmp(51388) := x"1000";
    tmp(51389) := x"0800";
    tmp(51390) := x"0800";
    tmp(51391) := x"0800";
    tmp(51392) := x"0800";
    tmp(51393) := x"0800";
    tmp(51394) := x"0800";
    tmp(51395) := x"0800";
    tmp(51396) := x"0800";
    tmp(51397) := x"1000";
    tmp(51398) := x"1000";
    tmp(51399) := x"1000";
    tmp(51400) := x"1000";
    tmp(51401) := x"1000";
    tmp(51402) := x"1000";
    tmp(51403) := x"0800";
    tmp(51404) := x"0800";
    tmp(51405) := x"0800";
    tmp(51406) := x"1000";
    tmp(51407) := x"1000";
    tmp(51408) := x"1000";
    tmp(51409) := x"1000";
    tmp(51410) := x"0800";
    tmp(51411) := x"0800";
    tmp(51412) := x"0800";
    tmp(51413) := x"0800";
    tmp(51414) := x"0800";
    tmp(51415) := x"1000";
    tmp(51416) := x"1000";
    tmp(51417) := x"1000";
    tmp(51418) := x"1000";
    tmp(51419) := x"1000";
    tmp(51420) := x"1000";
    tmp(51421) := x"1000";
    tmp(51422) := x"0800";
    tmp(51423) := x"0800";
    tmp(51424) := x"0800";
    tmp(51425) := x"0800";
    tmp(51426) := x"0800";
    tmp(51427) := x"0820";
    tmp(51428) := x"0820";
    tmp(51429) := x"0820";
    tmp(51430) := x"0800";
    tmp(51431) := x"1000";
    tmp(51432) := x"1000";
    tmp(51433) := x"1000";
    tmp(51434) := x"1800";
    tmp(51435) := x"1820";
    tmp(51436) := x"1820";
    tmp(51437) := x"1800";
    tmp(51438) := x"2020";
    tmp(51439) := x"3020";
    tmp(51440) := x"3820";
    tmp(51441) := x"3820";
    tmp(51442) := x"4020";
    tmp(51443) := x"3820";
    tmp(51444) := x"3000";
    tmp(51445) := x"2800";
    tmp(51446) := x"2000";
    tmp(51447) := x"2000";
    tmp(51448) := x"2820";
    tmp(51449) := x"4040";
    tmp(51450) := x"5841";
    tmp(51451) := x"5041";
    tmp(51452) := x"4841";
    tmp(51453) := x"4841";
    tmp(51454) := x"4020";
    tmp(51455) := x"4020";
    tmp(51456) := x"3020";
    tmp(51457) := x"3000";
    tmp(51458) := x"3000";
    tmp(51459) := x"3000";
    tmp(51460) := x"3800";
    tmp(51461) := x"4020";
    tmp(51462) := x"3820";
    tmp(51463) := x"3020";
    tmp(51464) := x"2820";
    tmp(51465) := x"2821";
    tmp(51466) := x"2021";
    tmp(51467) := x"1820";
    tmp(51468) := x"1000";
    tmp(51469) := x"1000";
    tmp(51470) := x"1000";
    tmp(51471) := x"0800";
    tmp(51472) := x"0000";
    tmp(51473) := x"0000";
    tmp(51474) := x"0000";
    tmp(51475) := x"0000";
    tmp(51476) := x"0000";
    tmp(51477) := x"0000";
    tmp(51478) := x"0000";
    tmp(51479) := x"0000";
    tmp(51480) := x"0000";
    tmp(51481) := x"0000";
    tmp(51482) := x"0000";
    tmp(51483) := x"0000";
    tmp(51484) := x"0000";
    tmp(51485) := x"0000";
    tmp(51486) := x"0000";
    tmp(51487) := x"0000";
    tmp(51488) := x"0000";
    tmp(51489) := x"0000";
    tmp(51490) := x"0000";
    tmp(51491) := x"0020";
    tmp(51492) := x"0020";
    tmp(51493) := x"0000";
    tmp(51494) := x"2882";
    tmp(51495) := x"b2ab";
    tmp(51496) := x"c30f";
    tmp(51497) := x"6946";
    tmp(51498) := x"89a7";
    tmp(51499) := x"cacc";
    tmp(51500) := x"8946";
    tmp(51501) := x"68c3";
    tmp(51502) := x"cb4e";
    tmp(51503) := x"922a";
    tmp(51504) := x"91e9";
    tmp(51505) := x"7105";
    tmp(51506) := x"8166";
    tmp(51507) := x"e390";
    tmp(51508) := x"4883";
    tmp(51509) := x"e30d";
    tmp(51510) := x"c2cd";
    tmp(51511) := x"91c8";
    tmp(51512) := x"50a3";
    tmp(51513) := x"9a8b";
    tmp(51514) := x"928c";
    tmp(51515) := x"92cd";
    tmp(51516) := x"722a";
    tmp(51517) := x"6a0a";
    tmp(51518) := x"59c8";
    tmp(51519) := x"5a09";
    tmp(51520) := x"728b";
    tmp(51521) := x"7a8b";
    tmp(51522) := x"5946";
    tmp(51523) := x"7166";
    tmp(51524) := x"ebf0";
    tmp(51525) := x"b1e9";
    tmp(51526) := x"2800";
    tmp(51527) := x"4000";
    tmp(51528) := x"5000";
    tmp(51529) := x"6800";
    tmp(51530) := x"6800";
    tmp(51531) := x"7000";
    tmp(51532) := x"6800";
    tmp(51533) := x"6800";
    tmp(51534) := x"8000";
    tmp(51535) := x"9000";
    tmp(51536) := x"9800";
    tmp(51537) := x"b020";
    tmp(51538) := x"a800";
    tmp(51539) := x"9800";
    tmp(51540) := x"a000";
    tmp(51541) := x"b820";
    tmp(51542) := x"b820";
    tmp(51543) := x"c820";
    tmp(51544) := x"b820";
    tmp(51545) := x"e040";
    tmp(51546) := x"f081";
    tmp(51547) := x"f8a1";
    tmp(51548) := x"5860";
    tmp(51549) := x"1020";
    tmp(51550) := x"0840";
    tmp(51551) := x"0840";
    tmp(51552) := x"0840";
    tmp(51553) := x"0840";
    tmp(51554) := x"0840";
    tmp(51555) := x"0840";
    tmp(51556) := x"0840";
    tmp(51557) := x"0840";
    tmp(51558) := x"0840";
    tmp(51559) := x"0840";
    tmp(51560) := x"0840";
    tmp(51561) := x"0840";
    tmp(51562) := x"0840";
    tmp(51563) := x"0840";
    tmp(51564) := x"0840";
    tmp(51565) := x"0840";
    tmp(51566) := x"0840";
    tmp(51567) := x"0840";
    tmp(51568) := x"0840";
    tmp(51569) := x"0840";
    tmp(51570) := x"0840";
    tmp(51571) := x"0840";
    tmp(51572) := x"0840";
    tmp(51573) := x"0840";
    tmp(51574) := x"0840";
    tmp(51575) := x"0840";
    tmp(51576) := x"0840";
    tmp(51577) := x"0840";
    tmp(51578) := x"0840";
    tmp(51579) := x"0840";
    tmp(51580) := x"0840";
    tmp(51581) := x"0840";
    tmp(51582) := x"0840";
    tmp(51583) := x"0840";
    tmp(51584) := x"0840";
    tmp(51585) := x"0840";
    tmp(51586) := x"0840";
    tmp(51587) := x"0840";
    tmp(51588) := x"0840";
    tmp(51589) := x"0840";
    tmp(51590) := x"0840";
    tmp(51591) := x"0840";
    tmp(51592) := x"0840";
    tmp(51593) := x"0840";
    tmp(51594) := x"0840";
    tmp(51595) := x"0840";
    tmp(51596) := x"0840";
    tmp(51597) := x"0840";
    tmp(51598) := x"0840";
    tmp(51599) := x"0840";
    tmp(51600) := x"0000";
    tmp(51601) := x"0860";
    tmp(51602) := x"0020";
    tmp(51603) := x"0000";
    tmp(51604) := x"0000";
    tmp(51605) := x"0000";
    tmp(51606) := x"0000";
    tmp(51607) := x"0000";
    tmp(51608) := x"0000";
    tmp(51609) := x"0000";
    tmp(51610) := x"0000";
    tmp(51611) := x"0820";
    tmp(51612) := x"0000";
    tmp(51613) := x"0000";
    tmp(51614) := x"0000";
    tmp(51615) := x"0000";
    tmp(51616) := x"0000";
    tmp(51617) := x"0000";
    tmp(51618) := x"0000";
    tmp(51619) := x"0800";
    tmp(51620) := x"0800";
    tmp(51621) := x"0800";
    tmp(51622) := x"0800";
    tmp(51623) := x"0800";
    tmp(51624) := x"0800";
    tmp(51625) := x"0800";
    tmp(51626) := x"0800";
    tmp(51627) := x"0800";
    tmp(51628) := x"0800";
    tmp(51629) := x"0800";
    tmp(51630) := x"0800";
    tmp(51631) := x"0800";
    tmp(51632) := x"0800";
    tmp(51633) := x"0800";
    tmp(51634) := x"0800";
    tmp(51635) := x"0800";
    tmp(51636) := x"0800";
    tmp(51637) := x"0800";
    tmp(51638) := x"0800";
    tmp(51639) := x"0800";
    tmp(51640) := x"1000";
    tmp(51641) := x"1000";
    tmp(51642) := x"0800";
    tmp(51643) := x"0800";
    tmp(51644) := x"0800";
    tmp(51645) := x"0800";
    tmp(51646) := x"1000";
    tmp(51647) := x"1800";
    tmp(51648) := x"2000";
    tmp(51649) := x"1800";
    tmp(51650) := x"1800";
    tmp(51651) := x"1800";
    tmp(51652) := x"1000";
    tmp(51653) := x"1000";
    tmp(51654) := x"1000";
    tmp(51655) := x"1000";
    tmp(51656) := x"1000";
    tmp(51657) := x"1000";
    tmp(51658) := x"1000";
    tmp(51659) := x"1000";
    tmp(51660) := x"1000";
    tmp(51661) := x"1000";
    tmp(51662) := x"1000";
    tmp(51663) := x"1000";
    tmp(51664) := x"1000";
    tmp(51665) := x"1000";
    tmp(51666) := x"1000";
    tmp(51667) := x"1020";
    tmp(51668) := x"1000";
    tmp(51669) := x"0800";
    tmp(51670) := x"1000";
    tmp(51671) := x"1800";
    tmp(51672) := x"2000";
    tmp(51673) := x"2000";
    tmp(51674) := x"2000";
    tmp(51675) := x"2800";
    tmp(51676) := x"2800";
    tmp(51677) := x"2000";
    tmp(51678) := x"2000";
    tmp(51679) := x"2800";
    tmp(51680) := x"2800";
    tmp(51681) := x"3020";
    tmp(51682) := x"3820";
    tmp(51683) := x"3020";
    tmp(51684) := x"3020";
    tmp(51685) := x"3020";
    tmp(51686) := x"2820";
    tmp(51687) := x"2820";
    tmp(51688) := x"2820";
    tmp(51689) := x"4841";
    tmp(51690) := x"5041";
    tmp(51691) := x"5041";
    tmp(51692) := x"5041";
    tmp(51693) := x"5041";
    tmp(51694) := x"4841";
    tmp(51695) := x"4041";
    tmp(51696) := x"3820";
    tmp(51697) := x"3020";
    tmp(51698) := x"3000";
    tmp(51699) := x"2800";
    tmp(51700) := x"2000";
    tmp(51701) := x"2800";
    tmp(51702) := x"3020";
    tmp(51703) := x"3020";
    tmp(51704) := x"2020";
    tmp(51705) := x"2020";
    tmp(51706) := x"1821";
    tmp(51707) := x"1820";
    tmp(51708) := x"1020";
    tmp(51709) := x"1000";
    tmp(51710) := x"0800";
    tmp(51711) := x"0800";
    tmp(51712) := x"0000";
    tmp(51713) := x"0000";
    tmp(51714) := x"0000";
    tmp(51715) := x"0000";
    tmp(51716) := x"0000";
    tmp(51717) := x"0000";
    tmp(51718) := x"0000";
    tmp(51719) := x"0000";
    tmp(51720) := x"0000";
    tmp(51721) := x"0000";
    tmp(51722) := x"0000";
    tmp(51723) := x"0000";
    tmp(51724) := x"0000";
    tmp(51725) := x"0000";
    tmp(51726) := x"0000";
    tmp(51727) := x"0000";
    tmp(51728) := x"0000";
    tmp(51729) := x"0000";
    tmp(51730) := x"0000";
    tmp(51731) := x"0020";
    tmp(51732) := x"0000";
    tmp(51733) := x"0820";
    tmp(51734) := x"b30c";
    tmp(51735) := x"d370";
    tmp(51736) := x"9a4b";
    tmp(51737) := x"7146";
    tmp(51738) := x"ca6a";
    tmp(51739) := x"4841";
    tmp(51740) := x"5061";
    tmp(51741) := x"b249";
    tmp(51742) := x"b2cd";
    tmp(51743) := x"6925";
    tmp(51744) := x"99e9";
    tmp(51745) := x"50a3";
    tmp(51746) := x"aa6a";
    tmp(51747) := x"fcf5";
    tmp(51748) := x"4062";
    tmp(51749) := x"eb4e";
    tmp(51750) := x"9a2a";
    tmp(51751) := x"99e8";
    tmp(51752) := x"40a3";
    tmp(51753) := x"a2ac";
    tmp(51754) := x"92ce";
    tmp(51755) := x"9330";
    tmp(51756) := x"51e9";
    tmp(51757) := x"3924";
    tmp(51758) := x"3923";
    tmp(51759) := x"3103";
    tmp(51760) := x"20a2";
    tmp(51761) := x"3104";
    tmp(51762) := x"6a2a";
    tmp(51763) := x"5105";
    tmp(51764) := x"a28b";
    tmp(51765) := x"f3f2";
    tmp(51766) := x"3000";
    tmp(51767) := x"3800";
    tmp(51768) := x"5000";
    tmp(51769) := x"6800";
    tmp(51770) := x"6800";
    tmp(51771) := x"7000";
    tmp(51772) := x"6800";
    tmp(51773) := x"6800";
    tmp(51774) := x"8800";
    tmp(51775) := x"a020";
    tmp(51776) := x"b020";
    tmp(51777) := x"c820";
    tmp(51778) := x"b020";
    tmp(51779) := x"9000";
    tmp(51780) := x"9800";
    tmp(51781) := x"b000";
    tmp(51782) := x"c020";
    tmp(51783) := x"d020";
    tmp(51784) := x"d020";
    tmp(51785) := x"e040";
    tmp(51786) := x"d840";
    tmp(51787) := x"e861";
    tmp(51788) := x"6061";
    tmp(51789) := x"1020";
    tmp(51790) := x"0840";
    tmp(51791) := x"0840";
    tmp(51792) := x"0840";
    tmp(51793) := x"0840";
    tmp(51794) := x"0840";
    tmp(51795) := x"0840";
    tmp(51796) := x"0840";
    tmp(51797) := x"0840";
    tmp(51798) := x"0840";
    tmp(51799) := x"0840";
    tmp(51800) := x"0840";
    tmp(51801) := x"0840";
    tmp(51802) := x"0840";
    tmp(51803) := x"0840";
    tmp(51804) := x"0840";
    tmp(51805) := x"0840";
    tmp(51806) := x"0840";
    tmp(51807) := x"0840";
    tmp(51808) := x"0840";
    tmp(51809) := x"0840";
    tmp(51810) := x"0840";
    tmp(51811) := x"0840";
    tmp(51812) := x"0840";
    tmp(51813) := x"0840";
    tmp(51814) := x"0840";
    tmp(51815) := x"0840";
    tmp(51816) := x"0840";
    tmp(51817) := x"0840";
    tmp(51818) := x"0840";
    tmp(51819) := x"0840";
    tmp(51820) := x"0840";
    tmp(51821) := x"0840";
    tmp(51822) := x"0840";
    tmp(51823) := x"0840";
    tmp(51824) := x"0840";
    tmp(51825) := x"0840";
    tmp(51826) := x"0840";
    tmp(51827) := x"0840";
    tmp(51828) := x"0840";
    tmp(51829) := x"0840";
    tmp(51830) := x"0840";
    tmp(51831) := x"0840";
    tmp(51832) := x"0840";
    tmp(51833) := x"0840";
    tmp(51834) := x"0840";
    tmp(51835) := x"0840";
    tmp(51836) := x"0840";
    tmp(51837) := x"0820";
    tmp(51838) := x"0820";
    tmp(51839) := x"0820";
    tmp(51840) := x"0000";
    tmp(51841) := x"0000";
    tmp(51842) := x"0000";
    tmp(51843) := x"0000";
    tmp(51844) := x"0000";
    tmp(51845) := x"0000";
    tmp(51846) := x"0000";
    tmp(51847) := x"0000";
    tmp(51848) := x"0000";
    tmp(51849) := x"0000";
    tmp(51850) := x"0000";
    tmp(51851) := x"0000";
    tmp(51852) := x"0000";
    tmp(51853) := x"0000";
    tmp(51854) := x"0000";
    tmp(51855) := x"0000";
    tmp(51856) := x"0800";
    tmp(51857) := x"0800";
    tmp(51858) := x"0800";
    tmp(51859) := x"0800";
    tmp(51860) := x"0800";
    tmp(51861) := x"0800";
    tmp(51862) := x"0800";
    tmp(51863) := x"0800";
    tmp(51864) := x"0800";
    tmp(51865) := x"0800";
    tmp(51866) := x"0800";
    tmp(51867) := x"0800";
    tmp(51868) := x"0800";
    tmp(51869) := x"0800";
    tmp(51870) := x"0800";
    tmp(51871) := x"0800";
    tmp(51872) := x"0800";
    tmp(51873) := x"0800";
    tmp(51874) := x"0800";
    tmp(51875) := x"0800";
    tmp(51876) := x"0800";
    tmp(51877) := x"0800";
    tmp(51878) := x"0800";
    tmp(51879) := x"0800";
    tmp(51880) := x"0800";
    tmp(51881) := x"0800";
    tmp(51882) := x"0800";
    tmp(51883) := x"0800";
    tmp(51884) := x"0800";
    tmp(51885) := x"1000";
    tmp(51886) := x"1800";
    tmp(51887) := x"2000";
    tmp(51888) := x"2000";
    tmp(51889) := x"2800";
    tmp(51890) := x"2800";
    tmp(51891) := x"2800";
    tmp(51892) := x"2800";
    tmp(51893) := x"2800";
    tmp(51894) := x"2800";
    tmp(51895) := x"2800";
    tmp(51896) := x"2000";
    tmp(51897) := x"2000";
    tmp(51898) := x"2000";
    tmp(51899) := x"2020";
    tmp(51900) := x"2000";
    tmp(51901) := x"2800";
    tmp(51902) := x"2000";
    tmp(51903) := x"2800";
    tmp(51904) := x"2800";
    tmp(51905) := x"2800";
    tmp(51906) := x"2800";
    tmp(51907) := x"3020";
    tmp(51908) := x"3020";
    tmp(51909) := x"2820";
    tmp(51910) := x"2000";
    tmp(51911) := x"2000";
    tmp(51912) := x"2000";
    tmp(51913) := x"2000";
    tmp(51914) := x"2800";
    tmp(51915) := x"2800";
    tmp(51916) := x"2800";
    tmp(51917) := x"2800";
    tmp(51918) := x"2000";
    tmp(51919) := x"2000";
    tmp(51920) := x"2000";
    tmp(51921) := x"2000";
    tmp(51922) := x"2800";
    tmp(51923) := x"2820";
    tmp(51924) := x"3020";
    tmp(51925) := x"3020";
    tmp(51926) := x"4041";
    tmp(51927) := x"3841";
    tmp(51928) := x"3820";
    tmp(51929) := x"4020";
    tmp(51930) := x"4020";
    tmp(51931) := x"4820";
    tmp(51932) := x"4841";
    tmp(51933) := x"4841";
    tmp(51934) := x"4041";
    tmp(51935) := x"4041";
    tmp(51936) := x"3821";
    tmp(51937) := x"3820";
    tmp(51938) := x"3820";
    tmp(51939) := x"3000";
    tmp(51940) := x"2000";
    tmp(51941) := x"1800";
    tmp(51942) := x"1800";
    tmp(51943) := x"2000";
    tmp(51944) := x"2820";
    tmp(51945) := x"1820";
    tmp(51946) := x"1020";
    tmp(51947) := x"1020";
    tmp(51948) := x"1020";
    tmp(51949) := x"0800";
    tmp(51950) := x"0800";
    tmp(51951) := x"0800";
    tmp(51952) := x"0000";
    tmp(51953) := x"0000";
    tmp(51954) := x"0000";
    tmp(51955) := x"0000";
    tmp(51956) := x"0000";
    tmp(51957) := x"0000";
    tmp(51958) := x"0000";
    tmp(51959) := x"0000";
    tmp(51960) := x"0000";
    tmp(51961) := x"0000";
    tmp(51962) := x"0000";
    tmp(51963) := x"0000";
    tmp(51964) := x"0000";
    tmp(51965) := x"0000";
    tmp(51966) := x"0000";
    tmp(51967) := x"0000";
    tmp(51968) := x"0000";
    tmp(51969) := x"0000";
    tmp(51970) := x"0000";
    tmp(51971) := x"0020";
    tmp(51972) := x"0000";
    tmp(51973) := x"5965";
    tmp(51974) := x"f454";
    tmp(51975) := x"b2ce";
    tmp(51976) := x"91c9";
    tmp(51977) := x"7925";
    tmp(51978) := x"a967";
    tmp(51979) := x"70a3";
    tmp(51980) := x"60a2";
    tmp(51981) := x"c2cc";
    tmp(51982) := x"9209";
    tmp(51983) := x"7987";
    tmp(51984) := x"dbb1";
    tmp(51985) := x"48a3";
    tmp(51986) := x"b26a";
    tmp(51987) := x"cacd";
    tmp(51988) := x"4062";
    tmp(51989) := x"fbf1";
    tmp(51990) := x"6946";
    tmp(51991) := x"8987";
    tmp(51992) := x"48a3";
    tmp(51993) := x"aaee";
    tmp(51994) := x"9b51";
    tmp(51995) := x"6a6c";
    tmp(51996) := x"4166";
    tmp(51997) := x"3103";
    tmp(51998) := x"28e2";
    tmp(51999) := x"18a2";
    tmp(52000) := x"18a2";
    tmp(52001) := x"1061";
    tmp(52002) := x"4186";
    tmp(52003) := x"7209";
    tmp(52004) := x"6146";
    tmp(52005) := x"ebb1";
    tmp(52006) := x"4841";
    tmp(52007) := x"3000";
    tmp(52008) := x"5000";
    tmp(52009) := x"6800";
    tmp(52010) := x"6800";
    tmp(52011) := x"7800";
    tmp(52012) := x"6800";
    tmp(52013) := x"6800";
    tmp(52014) := x"9000";
    tmp(52015) := x"a000";
    tmp(52016) := x"b020";
    tmp(52017) := x"c020";
    tmp(52018) := x"b020";
    tmp(52019) := x"9000";
    tmp(52020) := x"9800";
    tmp(52021) := x"b820";
    tmp(52022) := x"c020";
    tmp(52023) := x"c020";
    tmp(52024) := x"d820";
    tmp(52025) := x"e020";
    tmp(52026) := x"d020";
    tmp(52027) := x"e840";
    tmp(52028) := x"5840";
    tmp(52029) := x"1020";
    tmp(52030) := x"0820";
    tmp(52031) := x"0840";
    tmp(52032) := x"0840";
    tmp(52033) := x"0840";
    tmp(52034) := x"0840";
    tmp(52035) := x"0840";
    tmp(52036) := x"0840";
    tmp(52037) := x"0840";
    tmp(52038) := x"0840";
    tmp(52039) := x"0840";
    tmp(52040) := x"0840";
    tmp(52041) := x"0840";
    tmp(52042) := x"0840";
    tmp(52043) := x"0840";
    tmp(52044) := x"0840";
    tmp(52045) := x"0840";
    tmp(52046) := x"0840";
    tmp(52047) := x"0840";
    tmp(52048) := x"0840";
    tmp(52049) := x"0840";
    tmp(52050) := x"0840";
    tmp(52051) := x"0840";
    tmp(52052) := x"0840";
    tmp(52053) := x"0840";
    tmp(52054) := x"0840";
    tmp(52055) := x"0840";
    tmp(52056) := x"0840";
    tmp(52057) := x"0840";
    tmp(52058) := x"0840";
    tmp(52059) := x"0840";
    tmp(52060) := x"0840";
    tmp(52061) := x"0840";
    tmp(52062) := x"0840";
    tmp(52063) := x"0840";
    tmp(52064) := x"0840";
    tmp(52065) := x"0840";
    tmp(52066) := x"0840";
    tmp(52067) := x"0840";
    tmp(52068) := x"0840";
    tmp(52069) := x"0840";
    tmp(52070) := x"0840";
    tmp(52071) := x"0840";
    tmp(52072) := x"0840";
    tmp(52073) := x"0840";
    tmp(52074) := x"0840";
    tmp(52075) := x"0840";
    tmp(52076) := x"0820";
    tmp(52077) := x"0820";
    tmp(52078) := x"0820";
    tmp(52079) := x"0820";
    tmp(52080) := x"0000";
    tmp(52081) := x"0000";
    tmp(52082) := x"0000";
    tmp(52083) := x"0000";
    tmp(52084) := x"0000";
    tmp(52085) := x"0000";
    tmp(52086) := x"0000";
    tmp(52087) := x"0000";
    tmp(52088) := x"0000";
    tmp(52089) := x"0000";
    tmp(52090) := x"0000";
    tmp(52091) := x"0000";
    tmp(52092) := x"0000";
    tmp(52093) := x"0000";
    tmp(52094) := x"0800";
    tmp(52095) := x"0800";
    tmp(52096) := x"0820";
    tmp(52097) := x"0800";
    tmp(52098) := x"0800";
    tmp(52099) := x"1000";
    tmp(52100) := x"1000";
    tmp(52101) := x"1000";
    tmp(52102) := x"0800";
    tmp(52103) := x"0800";
    tmp(52104) := x"0800";
    tmp(52105) := x"0800";
    tmp(52106) := x"0800";
    tmp(52107) := x"0800";
    tmp(52108) := x"0800";
    tmp(52109) := x"0800";
    tmp(52110) := x"0800";
    tmp(52111) := x"0800";
    tmp(52112) := x"0800";
    tmp(52113) := x"0800";
    tmp(52114) := x"0800";
    tmp(52115) := x"0800";
    tmp(52116) := x"0800";
    tmp(52117) := x"0800";
    tmp(52118) := x"0800";
    tmp(52119) := x"0800";
    tmp(52120) := x"0800";
    tmp(52121) := x"0800";
    tmp(52122) := x"0800";
    tmp(52123) := x"1000";
    tmp(52124) := x"1000";
    tmp(52125) := x"1800";
    tmp(52126) := x"1800";
    tmp(52127) := x"1800";
    tmp(52128) := x"2000";
    tmp(52129) := x"2800";
    tmp(52130) := x"2800";
    tmp(52131) := x"3000";
    tmp(52132) := x"3000";
    tmp(52133) := x"3000";
    tmp(52134) := x"3000";
    tmp(52135) := x"3000";
    tmp(52136) := x"3000";
    tmp(52137) := x"3000";
    tmp(52138) := x"3000";
    tmp(52139) := x"3020";
    tmp(52140) := x"3000";
    tmp(52141) := x"3020";
    tmp(52142) := x"3820";
    tmp(52143) := x"3020";
    tmp(52144) := x"3000";
    tmp(52145) := x"3020";
    tmp(52146) := x"3020";
    tmp(52147) := x"3020";
    tmp(52148) := x"3020";
    tmp(52149) := x"3020";
    tmp(52150) := x"2800";
    tmp(52151) := x"2800";
    tmp(52152) := x"2000";
    tmp(52153) := x"2800";
    tmp(52154) := x"2800";
    tmp(52155) := x"2800";
    tmp(52156) := x"2800";
    tmp(52157) := x"2000";
    tmp(52158) := x"2000";
    tmp(52159) := x"1800";
    tmp(52160) := x"1800";
    tmp(52161) := x"1800";
    tmp(52162) := x"1800";
    tmp(52163) := x"1800";
    tmp(52164) := x"1000";
    tmp(52165) := x"1820";
    tmp(52166) := x"1020";
    tmp(52167) := x"1820";
    tmp(52168) := x"2020";
    tmp(52169) := x"3020";
    tmp(52170) := x"4020";
    tmp(52171) := x"4020";
    tmp(52172) := x"4020";
    tmp(52173) := x"4021";
    tmp(52174) := x"4041";
    tmp(52175) := x"3841";
    tmp(52176) := x"3021";
    tmp(52177) := x"3020";
    tmp(52178) := x"3820";
    tmp(52179) := x"3820";
    tmp(52180) := x"3000";
    tmp(52181) := x"2000";
    tmp(52182) := x"1000";
    tmp(52183) := x"1000";
    tmp(52184) := x"1800";
    tmp(52185) := x"2020";
    tmp(52186) := x"1000";
    tmp(52187) := x"1020";
    tmp(52188) := x"0800";
    tmp(52189) := x"0800";
    tmp(52190) := x"0800";
    tmp(52191) := x"0800";
    tmp(52192) := x"0000";
    tmp(52193) := x"0000";
    tmp(52194) := x"0000";
    tmp(52195) := x"0000";
    tmp(52196) := x"0000";
    tmp(52197) := x"0000";
    tmp(52198) := x"0000";
    tmp(52199) := x"0000";
    tmp(52200) := x"0000";
    tmp(52201) := x"0000";
    tmp(52202) := x"0000";
    tmp(52203) := x"0000";
    tmp(52204) := x"0000";
    tmp(52205) := x"0000";
    tmp(52206) := x"0000";
    tmp(52207) := x"0000";
    tmp(52208) := x"0000";
    tmp(52209) := x"0000";
    tmp(52210) := x"0000";
    tmp(52211) := x"0000";
    tmp(52212) := x"30a2";
    tmp(52213) := x"c32d";
    tmp(52214) := x"a26c";
    tmp(52215) := x"cb0f";
    tmp(52216) := x"50c4";
    tmp(52217) := x"c28b";
    tmp(52218) := x"e390";
    tmp(52219) := x"9187";
    tmp(52220) := x"8145";
    tmp(52221) := x"db0e";
    tmp(52222) := x"7125";
    tmp(52223) := x"91c8";
    tmp(52224) := x"aa6b";
    tmp(52225) := x"6905";
    tmp(52226) := x"dc52";
    tmp(52227) := x"c30e";
    tmp(52228) := x"4882";
    tmp(52229) := x"db70";
    tmp(52230) := x"48c3";
    tmp(52231) := x"99a7";
    tmp(52232) := x"48c3";
    tmp(52233) := x"bb71";
    tmp(52234) := x"82ae";
    tmp(52235) := x"4987";
    tmp(52236) := x"3924";
    tmp(52237) := x"2902";
    tmp(52238) := x"10a2";
    tmp(52239) := x"0841";
    tmp(52240) := x"0820";
    tmp(52241) := x"0841";
    tmp(52242) := x"1062";
    tmp(52243) := x"7acd";
    tmp(52244) := x"5967";
    tmp(52245) := x"a24b";
    tmp(52246) := x"70a3";
    tmp(52247) := x"3800";
    tmp(52248) := x"5800";
    tmp(52249) := x"6800";
    tmp(52250) := x"6800";
    tmp(52251) := x"8000";
    tmp(52252) := x"6800";
    tmp(52253) := x"7000";
    tmp(52254) := x"9020";
    tmp(52255) := x"a000";
    tmp(52256) := x"a000";
    tmp(52257) := x"c020";
    tmp(52258) := x"a000";
    tmp(52259) := x"a000";
    tmp(52260) := x"9800";
    tmp(52261) := x"b820";
    tmp(52262) := x"c820";
    tmp(52263) := x"c020";
    tmp(52264) := x"c820";
    tmp(52265) := x"d820";
    tmp(52266) := x"d020";
    tmp(52267) := x"e040";
    tmp(52268) := x"5040";
    tmp(52269) := x"0820";
    tmp(52270) := x"0840";
    tmp(52271) := x"0840";
    tmp(52272) := x"0840";
    tmp(52273) := x"0840";
    tmp(52274) := x"0840";
    tmp(52275) := x"0840";
    tmp(52276) := x"0840";
    tmp(52277) := x"0840";
    tmp(52278) := x"0840";
    tmp(52279) := x"0840";
    tmp(52280) := x"0840";
    tmp(52281) := x"0840";
    tmp(52282) := x"0820";
    tmp(52283) := x"0840";
    tmp(52284) := x"0840";
    tmp(52285) := x"0840";
    tmp(52286) := x"0840";
    tmp(52287) := x"0840";
    tmp(52288) := x"0840";
    tmp(52289) := x"0840";
    tmp(52290) := x"0840";
    tmp(52291) := x"0840";
    tmp(52292) := x"0840";
    tmp(52293) := x"0840";
    tmp(52294) := x"0840";
    tmp(52295) := x"0840";
    tmp(52296) := x"0840";
    tmp(52297) := x"0840";
    tmp(52298) := x"0840";
    tmp(52299) := x"0840";
    tmp(52300) := x"0840";
    tmp(52301) := x"0840";
    tmp(52302) := x"0840";
    tmp(52303) := x"0840";
    tmp(52304) := x"0840";
    tmp(52305) := x"0840";
    tmp(52306) := x"0840";
    tmp(52307) := x"0840";
    tmp(52308) := x"0840";
    tmp(52309) := x"0840";
    tmp(52310) := x"0840";
    tmp(52311) := x"0840";
    tmp(52312) := x"0840";
    tmp(52313) := x"0840";
    tmp(52314) := x"0840";
    tmp(52315) := x"0820";
    tmp(52316) := x"0820";
    tmp(52317) := x"0820";
    tmp(52318) := x"0820";
    tmp(52319) := x"0820";
    tmp(52320) := x"0000";
    tmp(52321) := x"0000";
    tmp(52322) := x"0000";
    tmp(52323) := x"0000";
    tmp(52324) := x"0000";
    tmp(52325) := x"0000";
    tmp(52326) := x"0000";
    tmp(52327) := x"0000";
    tmp(52328) := x"0000";
    tmp(52329) := x"0000";
    tmp(52330) := x"0000";
    tmp(52331) := x"0000";
    tmp(52332) := x"0000";
    tmp(52333) := x"0800";
    tmp(52334) := x"0800";
    tmp(52335) := x"0800";
    tmp(52336) := x"0800";
    tmp(52337) := x"0800";
    tmp(52338) := x"0800";
    tmp(52339) := x"1000";
    tmp(52340) := x"1000";
    tmp(52341) := x"1000";
    tmp(52342) := x"0800";
    tmp(52343) := x"0800";
    tmp(52344) := x"0800";
    tmp(52345) := x"0800";
    tmp(52346) := x"0800";
    tmp(52347) := x"0800";
    tmp(52348) := x"0800";
    tmp(52349) := x"0800";
    tmp(52350) := x"0800";
    tmp(52351) := x"0800";
    tmp(52352) := x"0800";
    tmp(52353) := x"0800";
    tmp(52354) := x"0800";
    tmp(52355) := x"0800";
    tmp(52356) := x"0800";
    tmp(52357) := x"0800";
    tmp(52358) := x"0800";
    tmp(52359) := x"0800";
    tmp(52360) := x"0800";
    tmp(52361) := x"1000";
    tmp(52362) := x"1800";
    tmp(52363) := x"1800";
    tmp(52364) := x"2000";
    tmp(52365) := x"2000";
    tmp(52366) := x"2000";
    tmp(52367) := x"2000";
    tmp(52368) := x"2000";
    tmp(52369) := x"2800";
    tmp(52370) := x"2800";
    tmp(52371) := x"2800";
    tmp(52372) := x"3000";
    tmp(52373) := x"3000";
    tmp(52374) := x"3000";
    tmp(52375) := x"3000";
    tmp(52376) := x"3000";
    tmp(52377) := x"3000";
    tmp(52378) := x"3820";
    tmp(52379) := x"3000";
    tmp(52380) := x"3000";
    tmp(52381) := x"3020";
    tmp(52382) := x"3020";
    tmp(52383) := x"3020";
    tmp(52384) := x"3020";
    tmp(52385) := x"3020";
    tmp(52386) := x"3020";
    tmp(52387) := x"3020";
    tmp(52388) := x"2820";
    tmp(52389) := x"2800";
    tmp(52390) := x"2800";
    tmp(52391) := x"2000";
    tmp(52392) := x"2000";
    tmp(52393) := x"2000";
    tmp(52394) := x"2000";
    tmp(52395) := x"2800";
    tmp(52396) := x"2000";
    tmp(52397) := x"2000";
    tmp(52398) := x"2000";
    tmp(52399) := x"1800";
    tmp(52400) := x"1800";
    tmp(52401) := x"1000";
    tmp(52402) := x"1000";
    tmp(52403) := x"1000";
    tmp(52404) := x"1020";
    tmp(52405) := x"1820";
    tmp(52406) := x"1820";
    tmp(52407) := x"2820";
    tmp(52408) := x"2820";
    tmp(52409) := x"2820";
    tmp(52410) := x"2820";
    tmp(52411) := x"3020";
    tmp(52412) := x"4021";
    tmp(52413) := x"4841";
    tmp(52414) := x"3841";
    tmp(52415) := x"3041";
    tmp(52416) := x"2841";
    tmp(52417) := x"2820";
    tmp(52418) := x"2820";
    tmp(52419) := x"3820";
    tmp(52420) := x"3800";
    tmp(52421) := x"3000";
    tmp(52422) := x"2820";
    tmp(52423) := x"1820";
    tmp(52424) := x"1000";
    tmp(52425) := x"0800";
    tmp(52426) := x"1000";
    tmp(52427) := x"1000";
    tmp(52428) := x"0800";
    tmp(52429) := x"0800";
    tmp(52430) := x"0800";
    tmp(52431) := x"0000";
    tmp(52432) := x"0000";
    tmp(52433) := x"0000";
    tmp(52434) := x"0000";
    tmp(52435) := x"0000";
    tmp(52436) := x"0000";
    tmp(52437) := x"0000";
    tmp(52438) := x"0000";
    tmp(52439) := x"0000";
    tmp(52440) := x"0000";
    tmp(52441) := x"0000";
    tmp(52442) := x"0000";
    tmp(52443) := x"0000";
    tmp(52444) := x"0000";
    tmp(52445) := x"0000";
    tmp(52446) := x"0000";
    tmp(52447) := x"0000";
    tmp(52448) := x"0000";
    tmp(52449) := x"0000";
    tmp(52450) := x"0000";
    tmp(52451) := x"2061";
    tmp(52452) := x"9a6a";
    tmp(52453) := x"bacd";
    tmp(52454) := x"c30e";
    tmp(52455) := x"91e9";
    tmp(52456) := x"7966";
    tmp(52457) := x"ebd1";
    tmp(52458) := x"cb4f";
    tmp(52459) := x"4882";
    tmp(52460) := x"e38f";
    tmp(52461) := x"aaac";
    tmp(52462) := x"8187";
    tmp(52463) := x"ebf2";
    tmp(52464) := x"48a3";
    tmp(52465) := x"8166";
    tmp(52466) := x"dbb1";
    tmp(52467) := x"db50";
    tmp(52468) := x"50a3";
    tmp(52469) := x"ec54";
    tmp(52470) := x"6925";
    tmp(52471) := x"a1c7";
    tmp(52472) := x"5904";
    tmp(52473) := x"c3f3";
    tmp(52474) := x"6a0b";
    tmp(52475) := x"51a7";
    tmp(52476) := x"3103";
    tmp(52477) := x"2102";
    tmp(52478) := x"0821";
    tmp(52479) := x"0000";
    tmp(52480) := x"0000";
    tmp(52481) := x"0821";
    tmp(52482) := x"0841";
    tmp(52483) := x"49c8";
    tmp(52484) := x"6a0b";
    tmp(52485) := x"6987";
    tmp(52486) := x"80e4";
    tmp(52487) := x"3800";
    tmp(52488) := x"5000";
    tmp(52489) := x"5800";
    tmp(52490) := x"7000";
    tmp(52491) := x"8820";
    tmp(52492) := x"6800";
    tmp(52493) := x"7000";
    tmp(52494) := x"9020";
    tmp(52495) := x"9800";
    tmp(52496) := x"a000";
    tmp(52497) := x"c020";
    tmp(52498) := x"a820";
    tmp(52499) := x"b020";
    tmp(52500) := x"b020";
    tmp(52501) := x"c020";
    tmp(52502) := x"c820";
    tmp(52503) := x"c020";
    tmp(52504) := x"c020";
    tmp(52505) := x"c820";
    tmp(52506) := x"d820";
    tmp(52507) := x"e041";
    tmp(52508) := x"4040";
    tmp(52509) := x"0820";
    tmp(52510) := x"0840";
    tmp(52511) := x"0840";
    tmp(52512) := x"0840";
    tmp(52513) := x"0840";
    tmp(52514) := x"0840";
    tmp(52515) := x"0840";
    tmp(52516) := x"0840";
    tmp(52517) := x"0840";
    tmp(52518) := x"0840";
    tmp(52519) := x"0840";
    tmp(52520) := x"0840";
    tmp(52521) := x"0840";
    tmp(52522) := x"0840";
    tmp(52523) := x"0840";
    tmp(52524) := x"0840";
    tmp(52525) := x"0840";
    tmp(52526) := x"0840";
    tmp(52527) := x"0840";
    tmp(52528) := x"0840";
    tmp(52529) := x"0840";
    tmp(52530) := x"0840";
    tmp(52531) := x"0840";
    tmp(52532) := x"0840";
    tmp(52533) := x"0840";
    tmp(52534) := x"0840";
    tmp(52535) := x"0840";
    tmp(52536) := x"0840";
    tmp(52537) := x"0840";
    tmp(52538) := x"0840";
    tmp(52539) := x"0840";
    tmp(52540) := x"0840";
    tmp(52541) := x"0840";
    tmp(52542) := x"0840";
    tmp(52543) := x"0840";
    tmp(52544) := x"0840";
    tmp(52545) := x"0840";
    tmp(52546) := x"0840";
    tmp(52547) := x"0840";
    tmp(52548) := x"0840";
    tmp(52549) := x"0840";
    tmp(52550) := x"0840";
    tmp(52551) := x"0840";
    tmp(52552) := x"0840";
    tmp(52553) := x"0820";
    tmp(52554) := x"0820";
    tmp(52555) := x"0820";
    tmp(52556) := x"0820";
    tmp(52557) := x"0820";
    tmp(52558) := x"0820";
    tmp(52559) := x"0820";
    tmp(52560) := x"0000";
    tmp(52561) := x"0000";
    tmp(52562) := x"0000";
    tmp(52563) := x"0000";
    tmp(52564) := x"0000";
    tmp(52565) := x"0000";
    tmp(52566) := x"0000";
    tmp(52567) := x"0000";
    tmp(52568) := x"0000";
    tmp(52569) := x"0000";
    tmp(52570) := x"0000";
    tmp(52571) := x"0800";
    tmp(52572) := x"0820";
    tmp(52573) := x"0800";
    tmp(52574) := x"0800";
    tmp(52575) := x"1000";
    tmp(52576) := x"1000";
    tmp(52577) := x"0800";
    tmp(52578) := x"1000";
    tmp(52579) := x"1000";
    tmp(52580) := x"0800";
    tmp(52581) := x"0800";
    tmp(52582) := x"0800";
    tmp(52583) := x"0800";
    tmp(52584) := x"0800";
    tmp(52585) := x"0800";
    tmp(52586) := x"0800";
    tmp(52587) := x"0800";
    tmp(52588) := x"0800";
    tmp(52589) := x"0800";
    tmp(52590) := x"0800";
    tmp(52591) := x"0800";
    tmp(52592) := x"0800";
    tmp(52593) := x"0800";
    tmp(52594) := x"0800";
    tmp(52595) := x"0800";
    tmp(52596) := x"0800";
    tmp(52597) := x"0800";
    tmp(52598) := x"0800";
    tmp(52599) := x"1000";
    tmp(52600) := x"1000";
    tmp(52601) := x"1800";
    tmp(52602) := x"2000";
    tmp(52603) := x"2000";
    tmp(52604) := x"2000";
    tmp(52605) := x"2000";
    tmp(52606) := x"2800";
    tmp(52607) := x"2800";
    tmp(52608) := x"2800";
    tmp(52609) := x"2800";
    tmp(52610) := x"3000";
    tmp(52611) := x"3000";
    tmp(52612) := x"3000";
    tmp(52613) := x"3000";
    tmp(52614) := x"3000";
    tmp(52615) := x"3000";
    tmp(52616) := x"3000";
    tmp(52617) := x"3000";
    tmp(52618) := x"3000";
    tmp(52619) := x"2800";
    tmp(52620) := x"3000";
    tmp(52621) := x"2800";
    tmp(52622) := x"3000";
    tmp(52623) := x"3020";
    tmp(52624) := x"3020";
    tmp(52625) := x"3020";
    tmp(52626) := x"3020";
    tmp(52627) := x"3020";
    tmp(52628) := x"2800";
    tmp(52629) := x"2000";
    tmp(52630) := x"2000";
    tmp(52631) := x"2000";
    tmp(52632) := x"2000";
    tmp(52633) := x"2000";
    tmp(52634) := x"2000";
    tmp(52635) := x"2000";
    tmp(52636) := x"2000";
    tmp(52637) := x"2000";
    tmp(52638) := x"2000";
    tmp(52639) := x"2000";
    tmp(52640) := x"1800";
    tmp(52641) := x"1800";
    tmp(52642) := x"1000";
    tmp(52643) := x"0800";
    tmp(52644) := x"1820";
    tmp(52645) := x"2820";
    tmp(52646) := x"3020";
    tmp(52647) := x"3020";
    tmp(52648) := x"3820";
    tmp(52649) := x"4020";
    tmp(52650) := x"4020";
    tmp(52651) := x"4821";
    tmp(52652) := x"4841";
    tmp(52653) := x"4841";
    tmp(52654) := x"4041";
    tmp(52655) := x"3841";
    tmp(52656) := x"3041";
    tmp(52657) := x"2861";
    tmp(52658) := x"2041";
    tmp(52659) := x"2020";
    tmp(52660) := x"3020";
    tmp(52661) := x"3000";
    tmp(52662) := x"3000";
    tmp(52663) := x"2820";
    tmp(52664) := x"1000";
    tmp(52665) := x"1020";
    tmp(52666) := x"0800";
    tmp(52667) := x"0800";
    tmp(52668) := x"0800";
    tmp(52669) := x"0800";
    tmp(52670) := x"0800";
    tmp(52671) := x"0000";
    tmp(52672) := x"0000";
    tmp(52673) := x"0000";
    tmp(52674) := x"0000";
    tmp(52675) := x"0000";
    tmp(52676) := x"0000";
    tmp(52677) := x"0000";
    tmp(52678) := x"0000";
    tmp(52679) := x"0000";
    tmp(52680) := x"0000";
    tmp(52681) := x"0000";
    tmp(52682) := x"0000";
    tmp(52683) := x"0000";
    tmp(52684) := x"0000";
    tmp(52685) := x"0000";
    tmp(52686) := x"0000";
    tmp(52687) := x"0000";
    tmp(52688) := x"0000";
    tmp(52689) := x"0000";
    tmp(52690) := x"0800";
    tmp(52691) := x"926a";
    tmp(52692) := x"c2ce";
    tmp(52693) := x"99ea";
    tmp(52694) := x"d30f";
    tmp(52695) := x"8187";
    tmp(52696) := x"b26b";
    tmp(52697) := x"ec13";
    tmp(52698) := x"aa6b";
    tmp(52699) := x"60e4";
    tmp(52700) := x"c2cd";
    tmp(52701) := x"8987";
    tmp(52702) := x"81a8";
    tmp(52703) := x"e391";
    tmp(52704) := x"5082";
    tmp(52705) := x"91a7";
    tmp(52706) := x"ebf2";
    tmp(52707) := x"8966";
    tmp(52708) := x"58a3";
    tmp(52709) := x"8125";
    tmp(52710) := x"4882";
    tmp(52711) := x"ba49";
    tmp(52712) := x"48a3";
    tmp(52713) := x"b371";
    tmp(52714) := x"6a0b";
    tmp(52715) := x"51a8";
    tmp(52716) := x"3123";
    tmp(52717) := x"2923";
    tmp(52718) := x"0841";
    tmp(52719) := x"0000";
    tmp(52720) := x"0000";
    tmp(52721) := x"0021";
    tmp(52722) := x"1062";
    tmp(52723) := x"3125";
    tmp(52724) := x"82ad";
    tmp(52725) := x"5105";
    tmp(52726) := x"4041";
    tmp(52727) := x"4800";
    tmp(52728) := x"6000";
    tmp(52729) := x"6000";
    tmp(52730) := x"7000";
    tmp(52731) := x"7000";
    tmp(52732) := x"6000";
    tmp(52733) := x"7000";
    tmp(52734) := x"a020";
    tmp(52735) := x"a000";
    tmp(52736) := x"a000";
    tmp(52737) := x"c820";
    tmp(52738) := x"b820";
    tmp(52739) := x"a820";
    tmp(52740) := x"c020";
    tmp(52741) := x"b820";
    tmp(52742) := x"c820";
    tmp(52743) := x"c820";
    tmp(52744) := x"c020";
    tmp(52745) := x"c820";
    tmp(52746) := x"e840";
    tmp(52747) := x"c861";
    tmp(52748) := x"2840";
    tmp(52749) := x"0820";
    tmp(52750) := x"0820";
    tmp(52751) := x"0820";
    tmp(52752) := x"0840";
    tmp(52753) := x"0840";
    tmp(52754) := x"0840";
    tmp(52755) := x"0840";
    tmp(52756) := x"0840";
    tmp(52757) := x"0840";
    tmp(52758) := x"0840";
    tmp(52759) := x"0840";
    tmp(52760) := x"0840";
    tmp(52761) := x"0840";
    tmp(52762) := x"0840";
    tmp(52763) := x"0840";
    tmp(52764) := x"0820";
    tmp(52765) := x"0840";
    tmp(52766) := x"0840";
    tmp(52767) := x"0840";
    tmp(52768) := x"0840";
    tmp(52769) := x"0840";
    tmp(52770) := x"0840";
    tmp(52771) := x"0840";
    tmp(52772) := x"0840";
    tmp(52773) := x"0840";
    tmp(52774) := x"0840";
    tmp(52775) := x"0840";
    tmp(52776) := x"0840";
    tmp(52777) := x"0840";
    tmp(52778) := x"0840";
    tmp(52779) := x"0840";
    tmp(52780) := x"0840";
    tmp(52781) := x"0840";
    tmp(52782) := x"0840";
    tmp(52783) := x"0840";
    tmp(52784) := x"0840";
    tmp(52785) := x"0840";
    tmp(52786) := x"0840";
    tmp(52787) := x"0840";
    tmp(52788) := x"0840";
    tmp(52789) := x"0840";
    tmp(52790) := x"0840";
    tmp(52791) := x"0840";
    tmp(52792) := x"0840";
    tmp(52793) := x"0820";
    tmp(52794) := x"0820";
    tmp(52795) := x"0820";
    tmp(52796) := x"0820";
    tmp(52797) := x"0820";
    tmp(52798) := x"0820";
    tmp(52799) := x"0820";
    tmp(52800) := x"0000";
    tmp(52801) := x"0000";
    tmp(52802) := x"0000";
    tmp(52803) := x"0000";
    tmp(52804) := x"0000";
    tmp(52805) := x"0000";
    tmp(52806) := x"0000";
    tmp(52807) := x"0000";
    tmp(52808) := x"0000";
    tmp(52809) := x"0800";
    tmp(52810) := x"0800";
    tmp(52811) := x"0800";
    tmp(52812) := x"0800";
    tmp(52813) := x"0800";
    tmp(52814) := x"0800";
    tmp(52815) := x"0800";
    tmp(52816) := x"1000";
    tmp(52817) := x"1000";
    tmp(52818) := x"1000";
    tmp(52819) := x"0800";
    tmp(52820) := x"0800";
    tmp(52821) := x"1000";
    tmp(52822) := x"1000";
    tmp(52823) := x"0800";
    tmp(52824) := x"0800";
    tmp(52825) := x"0800";
    tmp(52826) := x"0800";
    tmp(52827) := x"0800";
    tmp(52828) := x"0800";
    tmp(52829) := x"0800";
    tmp(52830) := x"0800";
    tmp(52831) := x"0800";
    tmp(52832) := x"0800";
    tmp(52833) := x"0800";
    tmp(52834) := x"0800";
    tmp(52835) := x"1000";
    tmp(52836) := x"1000";
    tmp(52837) := x"1000";
    tmp(52838) := x"1000";
    tmp(52839) := x"1800";
    tmp(52840) := x"2000";
    tmp(52841) := x"2000";
    tmp(52842) := x"2800";
    tmp(52843) := x"3020";
    tmp(52844) := x"3020";
    tmp(52845) := x"3020";
    tmp(52846) := x"3020";
    tmp(52847) := x"3020";
    tmp(52848) := x"2800";
    tmp(52849) := x"3000";
    tmp(52850) := x"3000";
    tmp(52851) := x"3000";
    tmp(52852) := x"3820";
    tmp(52853) := x"3820";
    tmp(52854) := x"3820";
    tmp(52855) := x"3820";
    tmp(52856) := x"3820";
    tmp(52857) := x"3800";
    tmp(52858) := x"3000";
    tmp(52859) := x"2800";
    tmp(52860) := x"2800";
    tmp(52861) := x"2800";
    tmp(52862) := x"3000";
    tmp(52863) := x"3000";
    tmp(52864) := x"3020";
    tmp(52865) := x"3020";
    tmp(52866) := x"3020";
    tmp(52867) := x"2800";
    tmp(52868) := x"2800";
    tmp(52869) := x"2800";
    tmp(52870) := x"2000";
    tmp(52871) := x"2000";
    tmp(52872) := x"2000";
    tmp(52873) := x"2000";
    tmp(52874) := x"2000";
    tmp(52875) := x"2000";
    tmp(52876) := x"2000";
    tmp(52877) := x"2000";
    tmp(52878) := x"2000";
    tmp(52879) := x"2000";
    tmp(52880) := x"1800";
    tmp(52881) := x"1800";
    tmp(52882) := x"1000";
    tmp(52883) := x"1820";
    tmp(52884) := x"2020";
    tmp(52885) := x"2020";
    tmp(52886) := x"2820";
    tmp(52887) := x"2820";
    tmp(52888) := x"2820";
    tmp(52889) := x"3020";
    tmp(52890) := x"3020";
    tmp(52891) := x"3020";
    tmp(52892) := x"3020";
    tmp(52893) := x"4841";
    tmp(52894) := x"4041";
    tmp(52895) := x"3841";
    tmp(52896) := x"3061";
    tmp(52897) := x"2861";
    tmp(52898) := x"2081";
    tmp(52899) := x"2882";
    tmp(52900) := x"2021";
    tmp(52901) := x"2020";
    tmp(52902) := x"2800";
    tmp(52903) := x"2820";
    tmp(52904) := x"1800";
    tmp(52905) := x"0800";
    tmp(52906) := x"0820";
    tmp(52907) := x"0800";
    tmp(52908) := x"0000";
    tmp(52909) := x"0800";
    tmp(52910) := x"0800";
    tmp(52911) := x"0000";
    tmp(52912) := x"0000";
    tmp(52913) := x"0000";
    tmp(52914) := x"0000";
    tmp(52915) := x"0000";
    tmp(52916) := x"0000";
    tmp(52917) := x"0000";
    tmp(52918) := x"0000";
    tmp(52919) := x"0000";
    tmp(52920) := x"0000";
    tmp(52921) := x"0000";
    tmp(52922) := x"0000";
    tmp(52923) := x"0000";
    tmp(52924) := x"0000";
    tmp(52925) := x"0000";
    tmp(52926) := x"0000";
    tmp(52927) := x"0000";
    tmp(52928) := x"0000";
    tmp(52929) := x"0000";
    tmp(52930) := x"5966";
    tmp(52931) := x"db91";
    tmp(52932) := x"89a8";
    tmp(52933) := x"db91";
    tmp(52934) := x"b24b";
    tmp(52935) := x"7946";
    tmp(52936) := x"ba8b";
    tmp(52937) := x"ec13";
    tmp(52938) := x"89a7";
    tmp(52939) := x"9a29";
    tmp(52940) := x"baac";
    tmp(52941) := x"60c4";
    tmp(52942) := x"c30d";
    tmp(52943) := x"8167";
    tmp(52944) := x"8125";
    tmp(52945) := x"e3d1";
    tmp(52946) := x"c24a";
    tmp(52947) := x"4041";
    tmp(52948) := x"ca08";
    tmp(52949) := x"5882";
    tmp(52950) := x"3861";
    tmp(52951) := x"8146";
    tmp(52952) := x"40a2";
    tmp(52953) := x"bb71";
    tmp(52954) := x"722c";
    tmp(52955) := x"4966";
    tmp(52956) := x"4144";
    tmp(52957) := x"3143";
    tmp(52958) := x"18a2";
    tmp(52959) := x"0841";
    tmp(52960) := x"0020";
    tmp(52961) := x"0861";
    tmp(52962) := x"1882";
    tmp(52963) := x"3105";
    tmp(52964) := x"722b";
    tmp(52965) := x"50a3";
    tmp(52966) := x"4020";
    tmp(52967) := x"5000";
    tmp(52968) := x"6000";
    tmp(52969) := x"5800";
    tmp(52970) := x"6800";
    tmp(52971) := x"7000";
    tmp(52972) := x"6000";
    tmp(52973) := x"7800";
    tmp(52974) := x"a020";
    tmp(52975) := x"9800";
    tmp(52976) := x"a000";
    tmp(52977) := x"c020";
    tmp(52978) := x"b820";
    tmp(52979) := x"a800";
    tmp(52980) := x"c820";
    tmp(52981) := x"c020";
    tmp(52982) := x"b820";
    tmp(52983) := x"c020";
    tmp(52984) := x"c820";
    tmp(52985) := x"e040";
    tmp(52986) := x"e840";
    tmp(52987) := x"c881";
    tmp(52988) := x"2840";
    tmp(52989) := x"0820";
    tmp(52990) := x"0820";
    tmp(52991) := x"0820";
    tmp(52992) := x"0840";
    tmp(52993) := x"0840";
    tmp(52994) := x"0840";
    tmp(52995) := x"0840";
    tmp(52996) := x"0840";
    tmp(52997) := x"0840";
    tmp(52998) := x"0840";
    tmp(52999) := x"0820";
    tmp(53000) := x"0840";
    tmp(53001) := x"0840";
    tmp(53002) := x"0840";
    tmp(53003) := x"0840";
    tmp(53004) := x"0840";
    tmp(53005) := x"0840";
    tmp(53006) := x"0840";
    tmp(53007) := x"0840";
    tmp(53008) := x"0840";
    tmp(53009) := x"0840";
    tmp(53010) := x"0840";
    tmp(53011) := x"0840";
    tmp(53012) := x"0840";
    tmp(53013) := x"0840";
    tmp(53014) := x"0840";
    tmp(53015) := x"0840";
    tmp(53016) := x"0840";
    tmp(53017) := x"0840";
    tmp(53018) := x"0840";
    tmp(53019) := x"0840";
    tmp(53020) := x"0840";
    tmp(53021) := x"0840";
    tmp(53022) := x"0840";
    tmp(53023) := x"0840";
    tmp(53024) := x"0840";
    tmp(53025) := x"0840";
    tmp(53026) := x"0840";
    tmp(53027) := x"0840";
    tmp(53028) := x"0820";
    tmp(53029) := x"0840";
    tmp(53030) := x"0820";
    tmp(53031) := x"0820";
    tmp(53032) := x"0820";
    tmp(53033) := x"0820";
    tmp(53034) := x"0820";
    tmp(53035) := x"0820";
    tmp(53036) := x"0820";
    tmp(53037) := x"0820";
    tmp(53038) := x"0820";
    tmp(53039) := x"0820";
    tmp(53040) := x"0000";
    tmp(53041) := x"0000";
    tmp(53042) := x"0000";
    tmp(53043) := x"0000";
    tmp(53044) := x"0000";
    tmp(53045) := x"0000";
    tmp(53046) := x"0000";
    tmp(53047) := x"0820";
    tmp(53048) := x"1021";
    tmp(53049) := x"0820";
    tmp(53050) := x"0800";
    tmp(53051) := x"0800";
    tmp(53052) := x"0800";
    tmp(53053) := x"0800";
    tmp(53054) := x"0800";
    tmp(53055) := x"1000";
    tmp(53056) := x"1000";
    tmp(53057) := x"1000";
    tmp(53058) := x"1000";
    tmp(53059) := x"1000";
    tmp(53060) := x"1000";
    tmp(53061) := x"1000";
    tmp(53062) := x"1000";
    tmp(53063) := x"1000";
    tmp(53064) := x"1000";
    tmp(53065) := x"1000";
    tmp(53066) := x"1000";
    tmp(53067) := x"0800";
    tmp(53068) := x"0800";
    tmp(53069) := x"0800";
    tmp(53070) := x"0800";
    tmp(53071) := x"1000";
    tmp(53072) := x"1000";
    tmp(53073) := x"1000";
    tmp(53074) := x"1000";
    tmp(53075) := x"1000";
    tmp(53076) := x"0800";
    tmp(53077) := x"0800";
    tmp(53078) := x"1000";
    tmp(53079) := x"1800";
    tmp(53080) := x"2000";
    tmp(53081) := x"2820";
    tmp(53082) := x"2820";
    tmp(53083) := x"3020";
    tmp(53084) := x"3020";
    tmp(53085) := x"3020";
    tmp(53086) := x"3020";
    tmp(53087) := x"3020";
    tmp(53088) := x"2800";
    tmp(53089) := x"3000";
    tmp(53090) := x"3000";
    tmp(53091) := x"3800";
    tmp(53092) := x"3820";
    tmp(53093) := x"4020";
    tmp(53094) := x"3820";
    tmp(53095) := x"3820";
    tmp(53096) := x"3800";
    tmp(53097) := x"3800";
    tmp(53098) := x"3000";
    tmp(53099) := x"3000";
    tmp(53100) := x"3000";
    tmp(53101) := x"2800";
    tmp(53102) := x"2800";
    tmp(53103) := x"3000";
    tmp(53104) := x"3000";
    tmp(53105) := x"2820";
    tmp(53106) := x"2820";
    tmp(53107) := x"2800";
    tmp(53108) := x"2800";
    tmp(53109) := x"2800";
    tmp(53110) := x"2800";
    tmp(53111) := x"2000";
    tmp(53112) := x"2000";
    tmp(53113) := x"2000";
    tmp(53114) := x"2000";
    tmp(53115) := x"2000";
    tmp(53116) := x"2000";
    tmp(53117) := x"2000";
    tmp(53118) := x"2000";
    tmp(53119) := x"1800";
    tmp(53120) := x"1800";
    tmp(53121) := x"1800";
    tmp(53122) := x"1000";
    tmp(53123) := x"1000";
    tmp(53124) := x"1800";
    tmp(53125) := x"2000";
    tmp(53126) := x"2000";
    tmp(53127) := x"2820";
    tmp(53128) := x"2800";
    tmp(53129) := x"2800";
    tmp(53130) := x"2820";
    tmp(53131) := x"2020";
    tmp(53132) := x"2020";
    tmp(53133) := x"2820";
    tmp(53134) := x"3020";
    tmp(53135) := x"3841";
    tmp(53136) := x"3041";
    tmp(53137) := x"2861";
    tmp(53138) := x"1861";
    tmp(53139) := x"1861";
    tmp(53140) := x"28a2";
    tmp(53141) := x"1841";
    tmp(53142) := x"1820";
    tmp(53143) := x"1800";
    tmp(53144) := x"1000";
    tmp(53145) := x"0800";
    tmp(53146) := x"0800";
    tmp(53147) := x"0820";
    tmp(53148) := x"0000";
    tmp(53149) := x"0000";
    tmp(53150) := x"0000";
    tmp(53151) := x"0000";
    tmp(53152) := x"0000";
    tmp(53153) := x"0000";
    tmp(53154) := x"0000";
    tmp(53155) := x"0000";
    tmp(53156) := x"0000";
    tmp(53157) := x"0000";
    tmp(53158) := x"0000";
    tmp(53159) := x"0000";
    tmp(53160) := x"0000";
    tmp(53161) := x"0000";
    tmp(53162) := x"0000";
    tmp(53163) := x"0000";
    tmp(53164) := x"0000";
    tmp(53165) := x"0000";
    tmp(53166) := x"0000";
    tmp(53167) := x"0000";
    tmp(53168) := x"0000";
    tmp(53169) := x"1041";
    tmp(53170) := x"bb0c";
    tmp(53171) := x"b26b";
    tmp(53172) := x"aa4b";
    tmp(53173) := x"db70";
    tmp(53174) := x"91e9";
    tmp(53175) := x"7126";
    tmp(53176) := x"aa4a";
    tmp(53177) := x"bacd";
    tmp(53178) := x"7125";
    tmp(53179) := x"8986";
    tmp(53180) := x"ba8b";
    tmp(53181) := x"68e4";
    tmp(53182) := x"fc33";
    tmp(53183) := x"6105";
    tmp(53184) := x"99a7";
    tmp(53185) := x"fdd9";
    tmp(53186) := x"8925";
    tmp(53187) := x"3820";
    tmp(53188) := x"9125";
    tmp(53189) := x"5062";
    tmp(53190) := x"60c3";
    tmp(53191) := x"99c7";
    tmp(53192) := x"4082";
    tmp(53193) := x"a2cd";
    tmp(53194) := x"92cf";
    tmp(53195) := x"5167";
    tmp(53196) := x"4986";
    tmp(53197) := x"3923";
    tmp(53198) := x"3123";
    tmp(53199) := x"18c2";
    tmp(53200) := x"18a2";
    tmp(53201) := x"18a2";
    tmp(53202) := x"20a2";
    tmp(53203) := x"3925";
    tmp(53204) := x"69a8";
    tmp(53205) := x"5061";
    tmp(53206) := x"4000";
    tmp(53207) := x"5000";
    tmp(53208) := x"5800";
    tmp(53209) := x"4800";
    tmp(53210) := x"6000";
    tmp(53211) := x"6800";
    tmp(53212) := x"6000";
    tmp(53213) := x"8800";
    tmp(53214) := x"9020";
    tmp(53215) := x"8800";
    tmp(53216) := x"9800";
    tmp(53217) := x"c020";
    tmp(53218) := x"b020";
    tmp(53219) := x"a800";
    tmp(53220) := x"c820";
    tmp(53221) := x"c820";
    tmp(53222) := x"c820";
    tmp(53223) := x"c020";
    tmp(53224) := x"c820";
    tmp(53225) := x"e040";
    tmp(53226) := x"f861";
    tmp(53227) := x"c081";
    tmp(53228) := x"2040";
    tmp(53229) := x"0820";
    tmp(53230) := x"0840";
    tmp(53231) := x"0820";
    tmp(53232) := x"0840";
    tmp(53233) := x"0840";
    tmp(53234) := x"0820";
    tmp(53235) := x"0840";
    tmp(53236) := x"0820";
    tmp(53237) := x"0840";
    tmp(53238) := x"0820";
    tmp(53239) := x"0840";
    tmp(53240) := x"0840";
    tmp(53241) := x"0840";
    tmp(53242) := x"0840";
    tmp(53243) := x"0820";
    tmp(53244) := x"0820";
    tmp(53245) := x"0840";
    tmp(53246) := x"0820";
    tmp(53247) := x"0840";
    tmp(53248) := x"0840";
    tmp(53249) := x"0840";
    tmp(53250) := x"0840";
    tmp(53251) := x"0840";
    tmp(53252) := x"0840";
    tmp(53253) := x"0840";
    tmp(53254) := x"0840";
    tmp(53255) := x"0840";
    tmp(53256) := x"0840";
    tmp(53257) := x"0840";
    tmp(53258) := x"0840";
    tmp(53259) := x"0840";
    tmp(53260) := x"0820";
    tmp(53261) := x"0840";
    tmp(53262) := x"0840";
    tmp(53263) := x"0840";
    tmp(53264) := x"0840";
    tmp(53265) := x"0840";
    tmp(53266) := x"0840";
    tmp(53267) := x"0840";
    tmp(53268) := x"0840";
    tmp(53269) := x"0840";
    tmp(53270) := x"0820";
    tmp(53271) := x"0820";
    tmp(53272) := x"0820";
    tmp(53273) := x"0820";
    tmp(53274) := x"0820";
    tmp(53275) := x"0820";
    tmp(53276) := x"0820";
    tmp(53277) := x"0820";
    tmp(53278) := x"0820";
    tmp(53279) := x"0820";
    tmp(53280) := x"0000";
    tmp(53281) := x"0000";
    tmp(53282) := x"0000";
    tmp(53283) := x"0000";
    tmp(53284) := x"0000";
    tmp(53285) := x"0800";
    tmp(53286) := x"0820";
    tmp(53287) := x"1020";
    tmp(53288) := x"0821";
    tmp(53289) := x"0820";
    tmp(53290) := x"0800";
    tmp(53291) := x"0800";
    tmp(53292) := x"0800";
    tmp(53293) := x"1000";
    tmp(53294) := x"1000";
    tmp(53295) := x"1000";
    tmp(53296) := x"1000";
    tmp(53297) := x"1000";
    tmp(53298) := x"1000";
    tmp(53299) := x"1000";
    tmp(53300) := x"1000";
    tmp(53301) := x"1000";
    tmp(53302) := x"1000";
    tmp(53303) := x"1000";
    tmp(53304) := x"1000";
    tmp(53305) := x"1000";
    tmp(53306) := x"1000";
    tmp(53307) := x"0800";
    tmp(53308) := x"0800";
    tmp(53309) := x"1000";
    tmp(53310) := x"1000";
    tmp(53311) := x"1000";
    tmp(53312) := x"1000";
    tmp(53313) := x"0800";
    tmp(53314) := x"0800";
    tmp(53315) := x"0800";
    tmp(53316) := x"0800";
    tmp(53317) := x"1000";
    tmp(53318) := x"1000";
    tmp(53319) := x"1800";
    tmp(53320) := x"1800";
    tmp(53321) := x"2000";
    tmp(53322) := x"2820";
    tmp(53323) := x"3020";
    tmp(53324) := x"3020";
    tmp(53325) := x"3820";
    tmp(53326) := x"3820";
    tmp(53327) := x"3820";
    tmp(53328) := x"3020";
    tmp(53329) := x"3000";
    tmp(53330) := x"3000";
    tmp(53331) := x"3000";
    tmp(53332) := x"3000";
    tmp(53333) := x"3000";
    tmp(53334) := x"3000";
    tmp(53335) := x"3000";
    tmp(53336) := x"3000";
    tmp(53337) := x"3000";
    tmp(53338) := x"3000";
    tmp(53339) := x"3800";
    tmp(53340) := x"3820";
    tmp(53341) := x"4020";
    tmp(53342) := x"4020";
    tmp(53343) := x"4020";
    tmp(53344) := x"3020";
    tmp(53345) := x"3000";
    tmp(53346) := x"3000";
    tmp(53347) := x"3000";
    tmp(53348) := x"2800";
    tmp(53349) := x"2800";
    tmp(53350) := x"2800";
    tmp(53351) := x"2000";
    tmp(53352) := x"2000";
    tmp(53353) := x"2000";
    tmp(53354) := x"2000";
    tmp(53355) := x"2000";
    tmp(53356) := x"2000";
    tmp(53357) := x"2000";
    tmp(53358) := x"2000";
    tmp(53359) := x"2000";
    tmp(53360) := x"2000";
    tmp(53361) := x"2000";
    tmp(53362) := x"1800";
    tmp(53363) := x"1800";
    tmp(53364) := x"2000";
    tmp(53365) := x"2000";
    tmp(53366) := x"2820";
    tmp(53367) := x"3020";
    tmp(53368) := x"3020";
    tmp(53369) := x"2800";
    tmp(53370) := x"2800";
    tmp(53371) := x"2020";
    tmp(53372) := x"1800";
    tmp(53373) := x"1000";
    tmp(53374) := x"1000";
    tmp(53375) := x"1800";
    tmp(53376) := x"1820";
    tmp(53377) := x"1820";
    tmp(53378) := x"1841";
    tmp(53379) := x"1041";
    tmp(53380) := x"1861";
    tmp(53381) := x"2082";
    tmp(53382) := x"1861";
    tmp(53383) := x"1841";
    tmp(53384) := x"0800";
    tmp(53385) := x"0800";
    tmp(53386) := x"0800";
    tmp(53387) := x"0000";
    tmp(53388) := x"0000";
    tmp(53389) := x"0000";
    tmp(53390) := x"0000";
    tmp(53391) := x"0000";
    tmp(53392) := x"0000";
    tmp(53393) := x"0000";
    tmp(53394) := x"0000";
    tmp(53395) := x"0000";
    tmp(53396) := x"0000";
    tmp(53397) := x"0000";
    tmp(53398) := x"0000";
    tmp(53399) := x"0000";
    tmp(53400) := x"0000";
    tmp(53401) := x"0000";
    tmp(53402) := x"0000";
    tmp(53403) := x"0000";
    tmp(53404) := x"0000";
    tmp(53405) := x"0000";
    tmp(53406) := x"0000";
    tmp(53407) := x"0000";
    tmp(53408) := x"0000";
    tmp(53409) := x"5966";
    tmp(53410) := x"caed";
    tmp(53411) := x"91a8";
    tmp(53412) := x"f3f2";
    tmp(53413) := x"aa2b";
    tmp(53414) := x"aa4c";
    tmp(53415) := x"89a8";
    tmp(53416) := x"a229";
    tmp(53417) := x"99a8";
    tmp(53418) := x"3041";
    tmp(53419) := x"ba08";
    tmp(53420) := x"b1c8";
    tmp(53421) := x"8125";
    tmp(53422) := x"eb0e";
    tmp(53423) := x"58a3";
    tmp(53424) := x"9187";
    tmp(53425) := x"fbf3";
    tmp(53426) := x"6882";
    tmp(53427) := x"5841";
    tmp(53428) := x"da2a";
    tmp(53429) := x"3020";
    tmp(53430) := x"70e3";
    tmp(53431) := x"99c8";
    tmp(53432) := x"2821";
    tmp(53433) := x"81a7";
    tmp(53434) := x"a2ef";
    tmp(53435) := x"69c9";
    tmp(53436) := x"5187";
    tmp(53437) := x"3924";
    tmp(53438) := x"4164";
    tmp(53439) := x"4984";
    tmp(53440) := x"4184";
    tmp(53441) := x"49a4";
    tmp(53442) := x"30c2";
    tmp(53443) := x"4946";
    tmp(53444) := x"6945";
    tmp(53445) := x"4020";
    tmp(53446) := x"4800";
    tmp(53447) := x"5800";
    tmp(53448) := x"5800";
    tmp(53449) := x"4800";
    tmp(53450) := x"6000";
    tmp(53451) := x"6800";
    tmp(53452) := x"6800";
    tmp(53453) := x"8800";
    tmp(53454) := x"8800";
    tmp(53455) := x"7800";
    tmp(53456) := x"9000";
    tmp(53457) := x"b020";
    tmp(53458) := x"b820";
    tmp(53459) := x"a820";
    tmp(53460) := x"c020";
    tmp(53461) := x"c820";
    tmp(53462) := x"e020";
    tmp(53463) := x"c820";
    tmp(53464) := x"c020";
    tmp(53465) := x"d820";
    tmp(53466) := x"e040";
    tmp(53467) := x"a840";
    tmp(53468) := x"2020";
    tmp(53469) := x"0820";
    tmp(53470) := x"0840";
    tmp(53471) := x"0820";
    tmp(53472) := x"0840";
    tmp(53473) := x"0820";
    tmp(53474) := x"0840";
    tmp(53475) := x"0840";
    tmp(53476) := x"0840";
    tmp(53477) := x"0840";
    tmp(53478) := x"0840";
    tmp(53479) := x"0840";
    tmp(53480) := x"0840";
    tmp(53481) := x"0840";
    tmp(53482) := x"0840";
    tmp(53483) := x"0820";
    tmp(53484) := x"0840";
    tmp(53485) := x"0840";
    tmp(53486) := x"0840";
    tmp(53487) := x"0840";
    tmp(53488) := x"0840";
    tmp(53489) := x"0840";
    tmp(53490) := x"0840";
    tmp(53491) := x"0840";
    tmp(53492) := x"0840";
    tmp(53493) := x"0840";
    tmp(53494) := x"0840";
    tmp(53495) := x"0840";
    tmp(53496) := x"0840";
    tmp(53497) := x"0840";
    tmp(53498) := x"0820";
    tmp(53499) := x"0820";
    tmp(53500) := x"0820";
    tmp(53501) := x"0840";
    tmp(53502) := x"0840";
    tmp(53503) := x"0840";
    tmp(53504) := x"0840";
    tmp(53505) := x"0840";
    tmp(53506) := x"0820";
    tmp(53507) := x"0820";
    tmp(53508) := x"0820";
    tmp(53509) := x"0820";
    tmp(53510) := x"0820";
    tmp(53511) := x"0820";
    tmp(53512) := x"0820";
    tmp(53513) := x"0820";
    tmp(53514) := x"0820";
    tmp(53515) := x"0820";
    tmp(53516) := x"0820";
    tmp(53517) := x"0820";
    tmp(53518) := x"0820";
    tmp(53519) := x"0820";
    tmp(53520) := x"0000";
    tmp(53521) := x"0000";
    tmp(53522) := x"0000";
    tmp(53523) := x"0000";
    tmp(53524) := x"0820";
    tmp(53525) := x"0820";
    tmp(53526) := x"0820";
    tmp(53527) := x"0820";
    tmp(53528) := x"0800";
    tmp(53529) := x"0800";
    tmp(53530) := x"0800";
    tmp(53531) := x"0800";
    tmp(53532) := x"1000";
    tmp(53533) := x"1000";
    tmp(53534) := x"1000";
    tmp(53535) := x"1000";
    tmp(53536) := x"1000";
    tmp(53537) := x"1000";
    tmp(53538) := x"1000";
    tmp(53539) := x"0800";
    tmp(53540) := x"0800";
    tmp(53541) := x"0800";
    tmp(53542) := x"0800";
    tmp(53543) := x"1000";
    tmp(53544) := x"1000";
    tmp(53545) := x"0800";
    tmp(53546) := x"0800";
    tmp(53547) := x"0800";
    tmp(53548) := x"0800";
    tmp(53549) := x"0800";
    tmp(53550) := x"0800";
    tmp(53551) := x"0800";
    tmp(53552) := x"0800";
    tmp(53553) := x"0800";
    tmp(53554) := x"1000";
    tmp(53555) := x"1000";
    tmp(53556) := x"1800";
    tmp(53557) := x"2000";
    tmp(53558) := x"2000";
    tmp(53559) := x"2000";
    tmp(53560) := x"1800";
    tmp(53561) := x"2000";
    tmp(53562) := x"2820";
    tmp(53563) := x"2820";
    tmp(53564) := x"2800";
    tmp(53565) := x"2800";
    tmp(53566) := x"2000";
    tmp(53567) := x"2000";
    tmp(53568) := x"2000";
    tmp(53569) := x"1800";
    tmp(53570) := x"2000";
    tmp(53571) := x"2000";
    tmp(53572) := x"2800";
    tmp(53573) := x"2800";
    tmp(53574) := x"2800";
    tmp(53575) := x"2800";
    tmp(53576) := x"2800";
    tmp(53577) := x"3000";
    tmp(53578) := x"3000";
    tmp(53579) := x"3000";
    tmp(53580) := x"3000";
    tmp(53581) := x"3000";
    tmp(53582) := x"3000";
    tmp(53583) := x"3000";
    tmp(53584) := x"3000";
    tmp(53585) := x"3000";
    tmp(53586) := x"3000";
    tmp(53587) := x"3000";
    tmp(53588) := x"2800";
    tmp(53589) := x"2800";
    tmp(53590) := x"2800";
    tmp(53591) := x"2800";
    tmp(53592) := x"2000";
    tmp(53593) := x"2800";
    tmp(53594) := x"2800";
    tmp(53595) := x"2800";
    tmp(53596) := x"2800";
    tmp(53597) := x"2800";
    tmp(53598) := x"2800";
    tmp(53599) := x"2000";
    tmp(53600) := x"2000";
    tmp(53601) := x"2000";
    tmp(53602) := x"2000";
    tmp(53603) := x"1800";
    tmp(53604) := x"2000";
    tmp(53605) := x"2000";
    tmp(53606) := x"2800";
    tmp(53607) := x"3020";
    tmp(53608) := x"3820";
    tmp(53609) := x"3820";
    tmp(53610) := x"3020";
    tmp(53611) := x"2800";
    tmp(53612) := x"2000";
    tmp(53613) := x"2020";
    tmp(53614) := x"2820";
    tmp(53615) := x"2820";
    tmp(53616) := x"2020";
    tmp(53617) := x"1800";
    tmp(53618) := x"1820";
    tmp(53619) := x"1020";
    tmp(53620) := x"1020";
    tmp(53621) := x"1841";
    tmp(53622) := x"2062";
    tmp(53623) := x"1841";
    tmp(53624) := x"1021";
    tmp(53625) := x"0800";
    tmp(53626) := x"0000";
    tmp(53627) := x"0000";
    tmp(53628) := x"0000";
    tmp(53629) := x"0000";
    tmp(53630) := x"0000";
    tmp(53631) := x"0000";
    tmp(53632) := x"0000";
    tmp(53633) := x"0000";
    tmp(53634) := x"0000";
    tmp(53635) := x"0000";
    tmp(53636) := x"0000";
    tmp(53637) := x"0000";
    tmp(53638) := x"0000";
    tmp(53639) := x"0000";
    tmp(53640) := x"0000";
    tmp(53641) := x"0000";
    tmp(53642) := x"0000";
    tmp(53643) := x"0000";
    tmp(53644) := x"0000";
    tmp(53645) := x"0000";
    tmp(53646) := x"0000";
    tmp(53647) := x"0000";
    tmp(53648) := x"1861";
    tmp(53649) := x"b2cb";
    tmp(53650) := x"ba6b";
    tmp(53651) := x"daed";
    tmp(53652) := x"d2ed";
    tmp(53653) := x"89a8";
    tmp(53654) := x"c2cd";
    tmp(53655) := x"7126";
    tmp(53656) := x"caed";
    tmp(53657) := x"60a3";
    tmp(53658) := x"4061";
    tmp(53659) := x"99a7";
    tmp(53660) := x"a9c7";
    tmp(53661) := x"70e4";
    tmp(53662) := x"c28b";
    tmp(53663) := x"58a3";
    tmp(53664) := x"99c8";
    tmp(53665) := x"fd7a";
    tmp(53666) := x"9125";
    tmp(53667) := x"70a3";
    tmp(53668) := x"f3d1";
    tmp(53669) := x"5062";
    tmp(53670) := x"4041";
    tmp(53671) := x"eb4d";
    tmp(53672) := x"5082";
    tmp(53673) := x"3862";
    tmp(53674) := x"aaad";
    tmp(53675) := x"a2ef";
    tmp(53676) := x"61a9";
    tmp(53677) := x"61e9";
    tmp(53678) := x"4986";
    tmp(53679) := x"3904";
    tmp(53680) := x"3924";
    tmp(53681) := x"3924";
    tmp(53682) := x"5186";
    tmp(53683) := x"69c8";
    tmp(53684) := x"60c3";
    tmp(53685) := x"2800";
    tmp(53686) := x"4800";
    tmp(53687) := x"5000";
    tmp(53688) := x"5000";
    tmp(53689) := x"5000";
    tmp(53690) := x"6000";
    tmp(53691) := x"6000";
    tmp(53692) := x"6800";
    tmp(53693) := x"7800";
    tmp(53694) := x"7800";
    tmp(53695) := x"8000";
    tmp(53696) := x"9000";
    tmp(53697) := x"a820";
    tmp(53698) := x"a800";
    tmp(53699) := x"b020";
    tmp(53700) := x"b000";
    tmp(53701) := x"c020";
    tmp(53702) := x"d020";
    tmp(53703) := x"d020";
    tmp(53704) := x"b820";
    tmp(53705) := x"d820";
    tmp(53706) := x"e040";
    tmp(53707) := x"a840";
    tmp(53708) := x"2020";
    tmp(53709) := x"0820";
    tmp(53710) := x"0840";
    tmp(53711) := x"0820";
    tmp(53712) := x"0840";
    tmp(53713) := x"0840";
    tmp(53714) := x"0840";
    tmp(53715) := x"0840";
    tmp(53716) := x"0840";
    tmp(53717) := x"0820";
    tmp(53718) := x"0840";
    tmp(53719) := x"0840";
    tmp(53720) := x"0820";
    tmp(53721) := x"0820";
    tmp(53722) := x"0820";
    tmp(53723) := x"0820";
    tmp(53724) := x"0840";
    tmp(53725) := x"0840";
    tmp(53726) := x"0840";
    tmp(53727) := x"0840";
    tmp(53728) := x"0820";
    tmp(53729) := x"0840";
    tmp(53730) := x"0840";
    tmp(53731) := x"0840";
    tmp(53732) := x"0820";
    tmp(53733) := x"0840";
    tmp(53734) := x"0840";
    tmp(53735) := x"0840";
    tmp(53736) := x"0840";
    tmp(53737) := x"0840";
    tmp(53738) := x"0820";
    tmp(53739) := x"0820";
    tmp(53740) := x"0820";
    tmp(53741) := x"0820";
    tmp(53742) := x"0820";
    tmp(53743) := x"0840";
    tmp(53744) := x"0820";
    tmp(53745) := x"0820";
    tmp(53746) := x"0820";
    tmp(53747) := x"0820";
    tmp(53748) := x"0820";
    tmp(53749) := x"0820";
    tmp(53750) := x"0820";
    tmp(53751) := x"0820";
    tmp(53752) := x"0820";
    tmp(53753) := x"0820";
    tmp(53754) := x"0820";
    tmp(53755) := x"0820";
    tmp(53756) := x"0820";
    tmp(53757) := x"0820";
    tmp(53758) := x"0820";
    tmp(53759) := x"0820";
    tmp(53760) := x"0000";
    tmp(53761) := x"0000";
    tmp(53762) := x"0800";
    tmp(53763) := x"0800";
    tmp(53764) := x"0800";
    tmp(53765) := x"0800";
    tmp(53766) := x"0800";
    tmp(53767) := x"0800";
    tmp(53768) := x"0800";
    tmp(53769) := x"0800";
    tmp(53770) := x"0800";
    tmp(53771) := x"0800";
    tmp(53772) := x"1000";
    tmp(53773) := x"0800";
    tmp(53774) := x"1000";
    tmp(53775) := x"1000";
    tmp(53776) := x"1000";
    tmp(53777) := x"1000";
    tmp(53778) := x"0800";
    tmp(53779) := x"0800";
    tmp(53780) := x"0800";
    tmp(53781) := x"0800";
    tmp(53782) := x"1000";
    tmp(53783) := x"0800";
    tmp(53784) := x"0800";
    tmp(53785) := x"0800";
    tmp(53786) := x"0800";
    tmp(53787) := x"0800";
    tmp(53788) := x"0800";
    tmp(53789) := x"0800";
    tmp(53790) := x"0800";
    tmp(53791) := x"0800";
    tmp(53792) := x"1000";
    tmp(53793) := x"1800";
    tmp(53794) := x"2000";
    tmp(53795) := x"2000";
    tmp(53796) := x"2000";
    tmp(53797) := x"2000";
    tmp(53798) := x"2000";
    tmp(53799) := x"2000";
    tmp(53800) := x"2000";
    tmp(53801) := x"2000";
    tmp(53802) := x"1800";
    tmp(53803) := x"1800";
    tmp(53804) := x"2000";
    tmp(53805) := x"2000";
    tmp(53806) := x"2000";
    tmp(53807) := x"2000";
    tmp(53808) := x"2800";
    tmp(53809) := x"2800";
    tmp(53810) := x"2800";
    tmp(53811) := x"2800";
    tmp(53812) := x"2800";
    tmp(53813) := x"2800";
    tmp(53814) := x"2800";
    tmp(53815) := x"2800";
    tmp(53816) := x"2800";
    tmp(53817) := x"3000";
    tmp(53818) := x"3000";
    tmp(53819) := x"3000";
    tmp(53820) := x"3000";
    tmp(53821) := x"3000";
    tmp(53822) := x"2800";
    tmp(53823) := x"2800";
    tmp(53824) := x"2800";
    tmp(53825) := x"2800";
    tmp(53826) := x"3000";
    tmp(53827) := x"2800";
    tmp(53828) := x"2800";
    tmp(53829) := x"2800";
    tmp(53830) := x"2800";
    tmp(53831) := x"2800";
    tmp(53832) := x"2800";
    tmp(53833) := x"2800";
    tmp(53834) := x"2800";
    tmp(53835) := x"2800";
    tmp(53836) := x"2800";
    tmp(53837) := x"2000";
    tmp(53838) := x"2000";
    tmp(53839) := x"2000";
    tmp(53840) := x"2000";
    tmp(53841) := x"2000";
    tmp(53842) := x"2000";
    tmp(53843) := x"1800";
    tmp(53844) := x"1800";
    tmp(53845) := x"1800";
    tmp(53846) := x"1800";
    tmp(53847) := x"2800";
    tmp(53848) := x"3020";
    tmp(53849) := x"3820";
    tmp(53850) := x"3820";
    tmp(53851) := x"2800";
    tmp(53852) := x"2000";
    tmp(53853) := x"3020";
    tmp(53854) := x"3020";
    tmp(53855) := x"3820";
    tmp(53856) := x"3020";
    tmp(53857) := x"2820";
    tmp(53858) := x"2000";
    tmp(53859) := x"1000";
    tmp(53860) := x"1000";
    tmp(53861) := x"1820";
    tmp(53862) := x"2020";
    tmp(53863) := x"2021";
    tmp(53864) := x"2021";
    tmp(53865) := x"1820";
    tmp(53866) := x"0800";
    tmp(53867) := x"0000";
    tmp(53868) := x"0000";
    tmp(53869) := x"0000";
    tmp(53870) := x"0000";
    tmp(53871) := x"0000";
    tmp(53872) := x"0000";
    tmp(53873) := x"0000";
    tmp(53874) := x"0000";
    tmp(53875) := x"0000";
    tmp(53876) := x"0000";
    tmp(53877) := x"0000";
    tmp(53878) := x"0000";
    tmp(53879) := x"0000";
    tmp(53880) := x"0000";
    tmp(53881) := x"0000";
    tmp(53882) := x"0000";
    tmp(53883) := x"0000";
    tmp(53884) := x"0000";
    tmp(53885) := x"0000";
    tmp(53886) := x"0000";
    tmp(53887) := x"1021";
    tmp(53888) := x"6985";
    tmp(53889) := x"91e8";
    tmp(53890) := x"c26b";
    tmp(53891) := x"db0e";
    tmp(53892) := x"aa2a";
    tmp(53893) := x"a22a";
    tmp(53894) := x"91c8";
    tmp(53895) := x"7946";
    tmp(53896) := x"caac";
    tmp(53897) := x"5082";
    tmp(53898) := x"68c3";
    tmp(53899) := x"f34d";
    tmp(53900) := x"9946";
    tmp(53901) := x"78c4";
    tmp(53902) := x"d28b";
    tmp(53903) := x"68a3";
    tmp(53904) := x"ba4a";
    tmp(53905) := x"fc14";
    tmp(53906) := x"a145";
    tmp(53907) := x"68a2";
    tmp(53908) := x"d30d";
    tmp(53909) := x"ca4a";
    tmp(53910) := x"2820";
    tmp(53911) := x"68c3";
    tmp(53912) := x"c24a";
    tmp(53913) := x"4862";
    tmp(53914) := x"6925";
    tmp(53915) := x"a28d";
    tmp(53916) := x"a2ef";
    tmp(53917) := x"7a4b";
    tmp(53918) := x"7a4b";
    tmp(53919) := x"61e9";
    tmp(53920) := x"6a2b";
    tmp(53921) := x"724b";
    tmp(53922) := x"722a";
    tmp(53923) := x"9209";
    tmp(53924) := x"3021";
    tmp(53925) := x"2800";
    tmp(53926) := x"4000";
    tmp(53927) := x"4800";
    tmp(53928) := x"4800";
    tmp(53929) := x"5000";
    tmp(53930) := x"6000";
    tmp(53931) := x"6800";
    tmp(53932) := x"6800";
    tmp(53933) := x"6800";
    tmp(53934) := x"7000";
    tmp(53935) := x"9000";
    tmp(53936) := x"8800";
    tmp(53937) := x"a000";
    tmp(53938) := x"a800";
    tmp(53939) := x"a000";
    tmp(53940) := x"a800";
    tmp(53941) := x"c020";
    tmp(53942) := x"c020";
    tmp(53943) := x"d820";
    tmp(53944) := x"c820";
    tmp(53945) := x"c820";
    tmp(53946) := x"e040";
    tmp(53947) := x"b861";
    tmp(53948) := x"2840";
    tmp(53949) := x"0820";
    tmp(53950) := x"0840";
    tmp(53951) := x"0840";
    tmp(53952) := x"0840";
    tmp(53953) := x"0840";
    tmp(53954) := x"0840";
    tmp(53955) := x"0820";
    tmp(53956) := x"0820";
    tmp(53957) := x"0820";
    tmp(53958) := x"0820";
    tmp(53959) := x"0820";
    tmp(53960) := x"0820";
    tmp(53961) := x"0820";
    tmp(53962) := x"0820";
    tmp(53963) := x"0820";
    tmp(53964) := x"0820";
    tmp(53965) := x"0840";
    tmp(53966) := x"0820";
    tmp(53967) := x"0820";
    tmp(53968) := x"0820";
    tmp(53969) := x"0820";
    tmp(53970) := x"0840";
    tmp(53971) := x"0820";
    tmp(53972) := x"0840";
    tmp(53973) := x"0820";
    tmp(53974) := x"0820";
    tmp(53975) := x"0820";
    tmp(53976) := x"0820";
    tmp(53977) := x"0820";
    tmp(53978) := x"0820";
    tmp(53979) := x"0820";
    tmp(53980) := x"0820";
    tmp(53981) := x"0820";
    tmp(53982) := x"0820";
    tmp(53983) := x"0820";
    tmp(53984) := x"0820";
    tmp(53985) := x"0820";
    tmp(53986) := x"0820";
    tmp(53987) := x"0820";
    tmp(53988) := x"0820";
    tmp(53989) := x"0820";
    tmp(53990) := x"0820";
    tmp(53991) := x"0820";
    tmp(53992) := x"0820";
    tmp(53993) := x"0820";
    tmp(53994) := x"0820";
    tmp(53995) := x"0820";
    tmp(53996) := x"0820";
    tmp(53997) := x"0820";
    tmp(53998) := x"0820";
    tmp(53999) := x"0820";
    tmp(54000) := x"0000";
    tmp(54001) := x"0820";
    tmp(54002) := x"0800";
    tmp(54003) := x"0000";
    tmp(54004) := x"0800";
    tmp(54005) := x"0800";
    tmp(54006) := x"0800";
    tmp(54007) := x"0800";
    tmp(54008) := x"0800";
    tmp(54009) := x"0800";
    tmp(54010) := x"0800";
    tmp(54011) := x"0800";
    tmp(54012) := x"0800";
    tmp(54013) := x"0800";
    tmp(54014) := x"0800";
    tmp(54015) := x"1000";
    tmp(54016) := x"0800";
    tmp(54017) := x"0800";
    tmp(54018) := x"0800";
    tmp(54019) := x"0800";
    tmp(54020) := x"0800";
    tmp(54021) := x"0800";
    tmp(54022) := x"1000";
    tmp(54023) := x"0800";
    tmp(54024) := x"0800";
    tmp(54025) := x"0800";
    tmp(54026) := x"0800";
    tmp(54027) := x"0800";
    tmp(54028) := x"0800";
    tmp(54029) := x"1000";
    tmp(54030) := x"1800";
    tmp(54031) := x"2000";
    tmp(54032) := x"2000";
    tmp(54033) := x"2000";
    tmp(54034) := x"2000";
    tmp(54035) := x"2000";
    tmp(54036) := x"2000";
    tmp(54037) := x"2000";
    tmp(54038) := x"2000";
    tmp(54039) := x"2000";
    tmp(54040) := x"2000";
    tmp(54041) := x"2000";
    tmp(54042) := x"2000";
    tmp(54043) := x"2000";
    tmp(54044) := x"2800";
    tmp(54045) := x"2800";
    tmp(54046) := x"2800";
    tmp(54047) := x"2800";
    tmp(54048) := x"2800";
    tmp(54049) := x"2800";
    tmp(54050) := x"2800";
    tmp(54051) := x"2800";
    tmp(54052) := x"2800";
    tmp(54053) := x"2800";
    tmp(54054) := x"2800";
    tmp(54055) := x"2800";
    tmp(54056) := x"2800";
    tmp(54057) := x"3000";
    tmp(54058) := x"2800";
    tmp(54059) := x"3000";
    tmp(54060) := x"3000";
    tmp(54061) := x"3000";
    tmp(54062) := x"2800";
    tmp(54063) := x"2800";
    tmp(54064) := x"2800";
    tmp(54065) := x"2800";
    tmp(54066) := x"2800";
    tmp(54067) := x"2800";
    tmp(54068) := x"2800";
    tmp(54069) := x"2800";
    tmp(54070) := x"2800";
    tmp(54071) := x"2800";
    tmp(54072) := x"2000";
    tmp(54073) := x"2000";
    tmp(54074) := x"2800";
    tmp(54075) := x"2800";
    tmp(54076) := x"2000";
    tmp(54077) := x"2000";
    tmp(54078) := x"2000";
    tmp(54079) := x"2000";
    tmp(54080) := x"2000";
    tmp(54081) := x"2000";
    tmp(54082) := x"2000";
    tmp(54083) := x"1800";
    tmp(54084) := x"1800";
    tmp(54085) := x"1000";
    tmp(54086) := x"1800";
    tmp(54087) := x"2000";
    tmp(54088) := x"3020";
    tmp(54089) := x"3820";
    tmp(54090) := x"3820";
    tmp(54091) := x"3020";
    tmp(54092) := x"2800";
    tmp(54093) := x"2820";
    tmp(54094) := x"3020";
    tmp(54095) := x"3020";
    tmp(54096) := x"3020";
    tmp(54097) := x"2820";
    tmp(54098) := x"2020";
    tmp(54099) := x"2020";
    tmp(54100) := x"2000";
    tmp(54101) := x"2000";
    tmp(54102) := x"2800";
    tmp(54103) := x"2000";
    tmp(54104) := x"2800";
    tmp(54105) := x"2820";
    tmp(54106) := x"2020";
    tmp(54107) := x"1000";
    tmp(54108) := x"0800";
    tmp(54109) := x"0000";
    tmp(54110) := x"0000";
    tmp(54111) := x"0000";
    tmp(54112) := x"0000";
    tmp(54113) := x"0000";
    tmp(54114) := x"0000";
    tmp(54115) := x"0000";
    tmp(54116) := x"0000";
    tmp(54117) := x"0000";
    tmp(54118) := x"0000";
    tmp(54119) := x"0000";
    tmp(54120) := x"0000";
    tmp(54121) := x"0000";
    tmp(54122) := x"0000";
    tmp(54123) := x"0000";
    tmp(54124) := x"0000";
    tmp(54125) := x"0000";
    tmp(54126) := x"0800";
    tmp(54127) := x"4904";
    tmp(54128) := x"9a29";
    tmp(54129) := x"99e8";
    tmp(54130) := x"c28c";
    tmp(54131) := x"db71";
    tmp(54132) := x"ba8d";
    tmp(54133) := x"99ea";
    tmp(54134) := x"8987";
    tmp(54135) := x"ba4b";
    tmp(54136) := x"b1e9";
    tmp(54137) := x"3841";
    tmp(54138) := x"58a2";
    tmp(54139) := x"d28b";
    tmp(54140) := x"9104";
    tmp(54141) := x"80e4";
    tmp(54142) := x"d229";
    tmp(54143) := x"5862";
    tmp(54144) := x"a1c8";
    tmp(54145) := x"eb90";
    tmp(54146) := x"78c3";
    tmp(54147) := x"4841";
    tmp(54148) := x"b1c7";
    tmp(54149) := x"68e4";
    tmp(54150) := x"b1c7";
    tmp(54151) := x"3021";
    tmp(54152) := x"99a7";
    tmp(54153) := x"a1c8";
    tmp(54154) := x"5083";
    tmp(54155) := x"50c4";
    tmp(54156) := x"aa6c";
    tmp(54157) := x"c391";
    tmp(54158) := x"92ee";
    tmp(54159) := x"826c";
    tmp(54160) := x"7a4b";
    tmp(54161) := x"71e9";
    tmp(54162) := x"8a4b";
    tmp(54163) := x"aa4a";
    tmp(54164) := x"2820";
    tmp(54165) := x"2800";
    tmp(54166) := x"3800";
    tmp(54167) := x"4000";
    tmp(54168) := x"4800";
    tmp(54169) := x"5800";
    tmp(54170) := x"6000";
    tmp(54171) := x"7000";
    tmp(54172) := x"7800";
    tmp(54173) := x"7000";
    tmp(54174) := x"7800";
    tmp(54175) := x"9000";
    tmp(54176) := x"8000";
    tmp(54177) := x"9000";
    tmp(54178) := x"a800";
    tmp(54179) := x"a000";
    tmp(54180) := x"a800";
    tmp(54181) := x"b820";
    tmp(54182) := x"c020";
    tmp(54183) := x"c820";
    tmp(54184) := x"d020";
    tmp(54185) := x"c020";
    tmp(54186) := x"d820";
    tmp(54187) := x"b040";
    tmp(54188) := x"2040";
    tmp(54189) := x"0820";
    tmp(54190) := x"0840";
    tmp(54191) := x"0820";
    tmp(54192) := x"0820";
    tmp(54193) := x"0820";
    tmp(54194) := x"0820";
    tmp(54195) := x"0820";
    tmp(54196) := x"0820";
    tmp(54197) := x"0820";
    tmp(54198) := x"0820";
    tmp(54199) := x"0820";
    tmp(54200) := x"0820";
    tmp(54201) := x"0820";
    tmp(54202) := x"0820";
    tmp(54203) := x"0840";
    tmp(54204) := x"0840";
    tmp(54205) := x"0840";
    tmp(54206) := x"0840";
    tmp(54207) := x"0840";
    tmp(54208) := x"0840";
    tmp(54209) := x"0840";
    tmp(54210) := x"0840";
    tmp(54211) := x"0840";
    tmp(54212) := x"0820";
    tmp(54213) := x"0820";
    tmp(54214) := x"0820";
    tmp(54215) := x"0820";
    tmp(54216) := x"0820";
    tmp(54217) := x"0820";
    tmp(54218) := x"0820";
    tmp(54219) := x"0820";
    tmp(54220) := x"0820";
    tmp(54221) := x"0820";
    tmp(54222) := x"0820";
    tmp(54223) := x"0820";
    tmp(54224) := x"0820";
    tmp(54225) := x"0820";
    tmp(54226) := x"0820";
    tmp(54227) := x"0820";
    tmp(54228) := x"0820";
    tmp(54229) := x"0820";
    tmp(54230) := x"0820";
    tmp(54231) := x"0820";
    tmp(54232) := x"0820";
    tmp(54233) := x"0820";
    tmp(54234) := x"0820";
    tmp(54235) := x"0820";
    tmp(54236) := x"0820";
    tmp(54237) := x"0820";
    tmp(54238) := x"0820";
    tmp(54239) := x"0820";
    tmp(54240) := x"0000";
    tmp(54241) := x"0000";
    tmp(54242) := x"0000";
    tmp(54243) := x"0000";
    tmp(54244) := x"0800";
    tmp(54245) := x"0800";
    tmp(54246) := x"0800";
    tmp(54247) := x"0800";
    tmp(54248) := x"0800";
    tmp(54249) := x"0800";
    tmp(54250) := x"0800";
    tmp(54251) := x"0800";
    tmp(54252) := x"0800";
    tmp(54253) := x"0800";
    tmp(54254) := x"0800";
    tmp(54255) := x"0800";
    tmp(54256) := x"0800";
    tmp(54257) := x"0800";
    tmp(54258) := x"0800";
    tmp(54259) := x"1000";
    tmp(54260) := x"1000";
    tmp(54261) := x"1000";
    tmp(54262) := x"1000";
    tmp(54263) := x"1000";
    tmp(54264) := x"1000";
    tmp(54265) := x"1000";
    tmp(54266) := x"1000";
    tmp(54267) := x"1000";
    tmp(54268) := x"1800";
    tmp(54269) := x"1800";
    tmp(54270) := x"1800";
    tmp(54271) := x"1800";
    tmp(54272) := x"1800";
    tmp(54273) := x"1800";
    tmp(54274) := x"1800";
    tmp(54275) := x"2000";
    tmp(54276) := x"2000";
    tmp(54277) := x"2000";
    tmp(54278) := x"2000";
    tmp(54279) := x"2000";
    tmp(54280) := x"2000";
    tmp(54281) := x"2000";
    tmp(54282) := x"2000";
    tmp(54283) := x"2800";
    tmp(54284) := x"2800";
    tmp(54285) := x"2800";
    tmp(54286) := x"3000";
    tmp(54287) := x"3000";
    tmp(54288) := x"2800";
    tmp(54289) := x"2800";
    tmp(54290) := x"2800";
    tmp(54291) := x"2800";
    tmp(54292) := x"2800";
    tmp(54293) := x"2800";
    tmp(54294) := x"2800";
    tmp(54295) := x"2800";
    tmp(54296) := x"3000";
    tmp(54297) := x"3000";
    tmp(54298) := x"3000";
    tmp(54299) := x"3000";
    tmp(54300) := x"3000";
    tmp(54301) := x"3000";
    tmp(54302) := x"3000";
    tmp(54303) := x"2800";
    tmp(54304) := x"2800";
    tmp(54305) := x"2000";
    tmp(54306) := x"2000";
    tmp(54307) := x"2000";
    tmp(54308) := x"2000";
    tmp(54309) := x"2000";
    tmp(54310) := x"2000";
    tmp(54311) := x"2000";
    tmp(54312) := x"2000";
    tmp(54313) := x"2000";
    tmp(54314) := x"2000";
    tmp(54315) := x"2000";
    tmp(54316) := x"2000";
    tmp(54317) := x"2000";
    tmp(54318) := x"2000";
    tmp(54319) := x"2000";
    tmp(54320) := x"2000";
    tmp(54321) := x"1800";
    tmp(54322) := x"1800";
    tmp(54323) := x"1800";
    tmp(54324) := x"1800";
    tmp(54325) := x"1000";
    tmp(54326) := x"1000";
    tmp(54327) := x"1000";
    tmp(54328) := x"1800";
    tmp(54329) := x"1800";
    tmp(54330) := x"2000";
    tmp(54331) := x"2000";
    tmp(54332) := x"1800";
    tmp(54333) := x"2000";
    tmp(54334) := x"2800";
    tmp(54335) := x"3000";
    tmp(54336) := x"3000";
    tmp(54337) := x"2820";
    tmp(54338) := x"2800";
    tmp(54339) := x"2000";
    tmp(54340) := x"2000";
    tmp(54341) := x"2000";
    tmp(54342) := x"2800";
    tmp(54343) := x"2800";
    tmp(54344) := x"2800";
    tmp(54345) := x"2800";
    tmp(54346) := x"2820";
    tmp(54347) := x"1820";
    tmp(54348) := x"0800";
    tmp(54349) := x"0800";
    tmp(54350) := x"0000";
    tmp(54351) := x"0000";
    tmp(54352) := x"0000";
    tmp(54353) := x"0000";
    tmp(54354) := x"0000";
    tmp(54355) := x"0000";
    tmp(54356) := x"0000";
    tmp(54357) := x"0000";
    tmp(54358) := x"0000";
    tmp(54359) := x"0000";
    tmp(54360) := x"0000";
    tmp(54361) := x"0000";
    tmp(54362) := x"0000";
    tmp(54363) := x"0000";
    tmp(54364) := x"0000";
    tmp(54365) := x"0000";
    tmp(54366) := x"2882";
    tmp(54367) := x"7186";
    tmp(54368) := x"8987";
    tmp(54369) := x"caac";
    tmp(54370) := x"c26c";
    tmp(54371) := x"db51";
    tmp(54372) := x"7968";
    tmp(54373) := x"b28c";
    tmp(54374) := x"ba4b";
    tmp(54375) := x"ba6b";
    tmp(54376) := x"ba09";
    tmp(54377) := x"3841";
    tmp(54378) := x"7904";
    tmp(54379) := x"b208";
    tmp(54380) := x"9104";
    tmp(54381) := x"9146";
    tmp(54382) := x"b9c8";
    tmp(54383) := x"4841";
    tmp(54384) := x"a9c8";
    tmp(54385) := x"a1e8";
    tmp(54386) := x"88c3";
    tmp(54387) := x"3820";
    tmp(54388) := x"e2eb";
    tmp(54389) := x"3841";
    tmp(54390) := x"c26a";
    tmp(54391) := x"99a7";
    tmp(54392) := x"4042";
    tmp(54393) := x"ca8c";
    tmp(54394) := x"9187";
    tmp(54395) := x"60c4";
    tmp(54396) := x"4062";
    tmp(54397) := x"7966";
    tmp(54398) := x"c36f";
    tmp(54399) := x"c391";
    tmp(54400) := x"a2cd";
    tmp(54401) := x"a28b";
    tmp(54402) := x"d38f";
    tmp(54403) := x"ba8a";
    tmp(54404) := x"2800";
    tmp(54405) := x"2000";
    tmp(54406) := x"3000";
    tmp(54407) := x"4000";
    tmp(54408) := x"4800";
    tmp(54409) := x"5000";
    tmp(54410) := x"6800";
    tmp(54411) := x"8820";
    tmp(54412) := x"7800";
    tmp(54413) := x"7800";
    tmp(54414) := x"8800";
    tmp(54415) := x"9020";
    tmp(54416) := x"8000";
    tmp(54417) := x"8800";
    tmp(54418) := x"a820";
    tmp(54419) := x"a000";
    tmp(54420) := x"b020";
    tmp(54421) := x"b820";
    tmp(54422) := x"b800";
    tmp(54423) := x"b820";
    tmp(54424) := x"c020";
    tmp(54425) := x"c820";
    tmp(54426) := x"d020";
    tmp(54427) := x"8840";
    tmp(54428) := x"1820";
    tmp(54429) := x"0820";
    tmp(54430) := x"0820";
    tmp(54431) := x"0820";
    tmp(54432) := x"0820";
    tmp(54433) := x"0820";
    tmp(54434) := x"0820";
    tmp(54435) := x"0820";
    tmp(54436) := x"0820";
    tmp(54437) := x"0820";
    tmp(54438) := x"0820";
    tmp(54439) := x"0820";
    tmp(54440) := x"0820";
    tmp(54441) := x"0820";
    tmp(54442) := x"0820";
    tmp(54443) := x"0840";
    tmp(54444) := x"0840";
    tmp(54445) := x"0840";
    tmp(54446) := x"0840";
    tmp(54447) := x"0840";
    tmp(54448) := x"0840";
    tmp(54449) := x"0840";
    tmp(54450) := x"0840";
    tmp(54451) := x"0840";
    tmp(54452) := x"0840";
    tmp(54453) := x"0820";
    tmp(54454) := x"0820";
    tmp(54455) := x"0820";
    tmp(54456) := x"0820";
    tmp(54457) := x"0820";
    tmp(54458) := x"0820";
    tmp(54459) := x"0820";
    tmp(54460) := x"0820";
    tmp(54461) := x"0820";
    tmp(54462) := x"0820";
    tmp(54463) := x"0820";
    tmp(54464) := x"0820";
    tmp(54465) := x"0820";
    tmp(54466) := x"0820";
    tmp(54467) := x"0820";
    tmp(54468) := x"0820";
    tmp(54469) := x"0820";
    tmp(54470) := x"0820";
    tmp(54471) := x"0820";
    tmp(54472) := x"0820";
    tmp(54473) := x"0820";
    tmp(54474) := x"0820";
    tmp(54475) := x"0820";
    tmp(54476) := x"0820";
    tmp(54477) := x"0820";
    tmp(54478) := x"0820";
    tmp(54479) := x"0820";
    tmp(54480) := x"0000";
    tmp(54481) := x"0000";
    tmp(54482) := x"0000";
    tmp(54483) := x"0800";
    tmp(54484) := x"0800";
    tmp(54485) := x"0800";
    tmp(54486) := x"0800";
    tmp(54487) := x"0800";
    tmp(54488) := x"0800";
    tmp(54489) := x"0800";
    tmp(54490) := x"0800";
    tmp(54491) := x"0800";
    tmp(54492) := x"0800";
    tmp(54493) := x"0800";
    tmp(54494) := x"0800";
    tmp(54495) := x"1000";
    tmp(54496) := x"1000";
    tmp(54497) := x"1000";
    tmp(54498) := x"1000";
    tmp(54499) := x"1000";
    tmp(54500) := x"1000";
    tmp(54501) := x"1000";
    tmp(54502) := x"1000";
    tmp(54503) := x"1000";
    tmp(54504) := x"1000";
    tmp(54505) := x"1800";
    tmp(54506) := x"1800";
    tmp(54507) := x"1800";
    tmp(54508) := x"1800";
    tmp(54509) := x"1800";
    tmp(54510) := x"1800";
    tmp(54511) := x"1800";
    tmp(54512) := x"1800";
    tmp(54513) := x"1800";
    tmp(54514) := x"1800";
    tmp(54515) := x"2000";
    tmp(54516) := x"2000";
    tmp(54517) := x"2000";
    tmp(54518) := x"2000";
    tmp(54519) := x"2000";
    tmp(54520) := x"2800";
    tmp(54521) := x"2800";
    tmp(54522) := x"2800";
    tmp(54523) := x"3000";
    tmp(54524) := x"3000";
    tmp(54525) := x"3000";
    tmp(54526) := x"3000";
    tmp(54527) := x"2800";
    tmp(54528) := x"2800";
    tmp(54529) := x"2800";
    tmp(54530) := x"2800";
    tmp(54531) := x"2800";
    tmp(54532) := x"2800";
    tmp(54533) := x"2800";
    tmp(54534) := x"2800";
    tmp(54535) := x"2800";
    tmp(54536) := x"3000";
    tmp(54537) := x"3000";
    tmp(54538) := x"3000";
    tmp(54539) := x"3000";
    tmp(54540) := x"3800";
    tmp(54541) := x"3800";
    tmp(54542) := x"3800";
    tmp(54543) := x"3000";
    tmp(54544) := x"3000";
    tmp(54545) := x"2800";
    tmp(54546) := x"2000";
    tmp(54547) := x"2000";
    tmp(54548) := x"2000";
    tmp(54549) := x"2000";
    tmp(54550) := x"1800";
    tmp(54551) := x"2000";
    tmp(54552) := x"2000";
    tmp(54553) := x"2000";
    tmp(54554) := x"2000";
    tmp(54555) := x"2000";
    tmp(54556) := x"1800";
    tmp(54557) := x"1800";
    tmp(54558) := x"1800";
    tmp(54559) := x"1800";
    tmp(54560) := x"1800";
    tmp(54561) := x"1800";
    tmp(54562) := x"1800";
    tmp(54563) := x"1800";
    tmp(54564) := x"1800";
    tmp(54565) := x"1800";
    tmp(54566) := x"1000";
    tmp(54567) := x"0800";
    tmp(54568) := x"0800";
    tmp(54569) := x"0800";
    tmp(54570) := x"0800";
    tmp(54571) := x"0800";
    tmp(54572) := x"0800";
    tmp(54573) := x"0800";
    tmp(54574) := x"1000";
    tmp(54575) := x"2000";
    tmp(54576) := x"2800";
    tmp(54577) := x"3000";
    tmp(54578) := x"2800";
    tmp(54579) := x"2000";
    tmp(54580) := x"2000";
    tmp(54581) := x"2000";
    tmp(54582) := x"1800";
    tmp(54583) := x"2000";
    tmp(54584) := x"2000";
    tmp(54585) := x"1800";
    tmp(54586) := x"1000";
    tmp(54587) := x"1000";
    tmp(54588) := x"0800";
    tmp(54589) := x"0800";
    tmp(54590) := x"0800";
    tmp(54591) := x"0800";
    tmp(54592) := x"0000";
    tmp(54593) := x"0000";
    tmp(54594) := x"0000";
    tmp(54595) := x"0000";
    tmp(54596) := x"0000";
    tmp(54597) := x"0000";
    tmp(54598) := x"0000";
    tmp(54599) := x"0000";
    tmp(54600) := x"0000";
    tmp(54601) := x"0000";
    tmp(54602) := x"0000";
    tmp(54603) := x"0000";
    tmp(54604) := x"0000";
    tmp(54605) := x"2081";
    tmp(54606) := x"5944";
    tmp(54607) := x"6945";
    tmp(54608) := x"99e8";
    tmp(54609) := x"d2ce";
    tmp(54610) := x"ca8d";
    tmp(54611) := x"8988";
    tmp(54612) := x"91a8";
    tmp(54613) := x"ebf2";
    tmp(54614) := x"a20a";
    tmp(54615) := x"c2cc";
    tmp(54616) := x"70e4";
    tmp(54617) := x"3021";
    tmp(54618) := x"e32d";
    tmp(54619) := x"ebd1";
    tmp(54620) := x"b22a";
    tmp(54621) := x"a9e9";
    tmp(54622) := x"9146";
    tmp(54623) := x"5041";
    tmp(54624) := x"cacc";
    tmp(54625) := x"a1e8";
    tmp(54626) := x"6882";
    tmp(54627) := x"3820";
    tmp(54628) := x"daec";
    tmp(54629) := x"8966";
    tmp(54630) := x"4042";
    tmp(54631) := x"fcd5";
    tmp(54632) := x"68c4";
    tmp(54633) := x"68a3";
    tmp(54634) := x"9126";
    tmp(54635) := x"7904";
    tmp(54636) := x"5061";
    tmp(54637) := x"2820";
    tmp(54638) := x"7104";
    tmp(54639) := x"baec";
    tmp(54640) := x"d390";
    tmp(54641) := x"cb4e";
    tmp(54642) := x"c32d";
    tmp(54643) := x"a1e7";
    tmp(54644) := x"2000";
    tmp(54645) := x"2000";
    tmp(54646) := x"3000";
    tmp(54647) := x"3800";
    tmp(54648) := x"4000";
    tmp(54649) := x"5000";
    tmp(54650) := x"7800";
    tmp(54651) := x"8800";
    tmp(54652) := x"7000";
    tmp(54653) := x"8000";
    tmp(54654) := x"9020";
    tmp(54655) := x"9820";
    tmp(54656) := x"8800";
    tmp(54657) := x"8000";
    tmp(54658) := x"a820";
    tmp(54659) := x"a820";
    tmp(54660) := x"c020";
    tmp(54661) := x"b820";
    tmp(54662) := x"b820";
    tmp(54663) := x"b820";
    tmp(54664) := x"b800";
    tmp(54665) := x"c020";
    tmp(54666) := x"c020";
    tmp(54667) := x"7040";
    tmp(54668) := x"1020";
    tmp(54669) := x"0820";
    tmp(54670) := x"0820";
    tmp(54671) := x"0820";
    tmp(54672) := x"0820";
    tmp(54673) := x"0820";
    tmp(54674) := x"0820";
    tmp(54675) := x"0820";
    tmp(54676) := x"0820";
    tmp(54677) := x"0820";
    tmp(54678) := x"0820";
    tmp(54679) := x"0820";
    tmp(54680) := x"0820";
    tmp(54681) := x"0820";
    tmp(54682) := x"0840";
    tmp(54683) := x"0840";
    tmp(54684) := x"0840";
    tmp(54685) := x"0840";
    tmp(54686) := x"0840";
    tmp(54687) := x"0840";
    tmp(54688) := x"0840";
    tmp(54689) := x"0840";
    tmp(54690) := x"0840";
    tmp(54691) := x"0840";
    tmp(54692) := x"0840";
    tmp(54693) := x"0820";
    tmp(54694) := x"0820";
    tmp(54695) := x"0820";
    tmp(54696) := x"0820";
    tmp(54697) := x"0820";
    tmp(54698) := x"0820";
    tmp(54699) := x"0820";
    tmp(54700) := x"0820";
    tmp(54701) := x"0820";
    tmp(54702) := x"0820";
    tmp(54703) := x"0820";
    tmp(54704) := x"0820";
    tmp(54705) := x"0820";
    tmp(54706) := x"0820";
    tmp(54707) := x"0820";
    tmp(54708) := x"0820";
    tmp(54709) := x"0820";
    tmp(54710) := x"0820";
    tmp(54711) := x"0820";
    tmp(54712) := x"0820";
    tmp(54713) := x"0820";
    tmp(54714) := x"0820";
    tmp(54715) := x"0820";
    tmp(54716) := x"0820";
    tmp(54717) := x"0820";
    tmp(54718) := x"0820";
    tmp(54719) := x"0820";
    tmp(54720) := x"0000";
    tmp(54721) := x"0000";
    tmp(54722) := x"0000";
    tmp(54723) := x"0800";
    tmp(54724) := x"0000";
    tmp(54725) := x"0800";
    tmp(54726) := x"0800";
    tmp(54727) := x"0800";
    tmp(54728) := x"0800";
    tmp(54729) := x"0800";
    tmp(54730) := x"0800";
    tmp(54731) := x"0800";
    tmp(54732) := x"1000";
    tmp(54733) := x"1000";
    tmp(54734) := x"1000";
    tmp(54735) := x"1800";
    tmp(54736) := x"1800";
    tmp(54737) := x"1000";
    tmp(54738) := x"1000";
    tmp(54739) := x"1000";
    tmp(54740) := x"1800";
    tmp(54741) := x"1800";
    tmp(54742) := x"1800";
    tmp(54743) := x"1800";
    tmp(54744) := x"1800";
    tmp(54745) := x"1800";
    tmp(54746) := x"2000";
    tmp(54747) := x"2000";
    tmp(54748) := x"1800";
    tmp(54749) := x"1800";
    tmp(54750) := x"1800";
    tmp(54751) := x"1800";
    tmp(54752) := x"1800";
    tmp(54753) := x"2000";
    tmp(54754) := x"2000";
    tmp(54755) := x"2000";
    tmp(54756) := x"2000";
    tmp(54757) := x"2000";
    tmp(54758) := x"2000";
    tmp(54759) := x"2800";
    tmp(54760) := x"2800";
    tmp(54761) := x"3000";
    tmp(54762) := x"3000";
    tmp(54763) := x"3000";
    tmp(54764) := x"3000";
    tmp(54765) := x"3000";
    tmp(54766) := x"2800";
    tmp(54767) := x"2800";
    tmp(54768) := x"2800";
    tmp(54769) := x"2800";
    tmp(54770) := x"2800";
    tmp(54771) := x"2800";
    tmp(54772) := x"2800";
    tmp(54773) := x"2800";
    tmp(54774) := x"2800";
    tmp(54775) := x"2800";
    tmp(54776) := x"2800";
    tmp(54777) := x"3000";
    tmp(54778) := x"3000";
    tmp(54779) := x"3000";
    tmp(54780) := x"3800";
    tmp(54781) := x"3000";
    tmp(54782) := x"3800";
    tmp(54783) := x"3000";
    tmp(54784) := x"2800";
    tmp(54785) := x"2800";
    tmp(54786) := x"2800";
    tmp(54787) := x"2000";
    tmp(54788) := x"2000";
    tmp(54789) := x"1800";
    tmp(54790) := x"1800";
    tmp(54791) := x"1800";
    tmp(54792) := x"1800";
    tmp(54793) := x"1800";
    tmp(54794) := x"2000";
    tmp(54795) := x"1800";
    tmp(54796) := x"1800";
    tmp(54797) := x"1800";
    tmp(54798) := x"1800";
    tmp(54799) := x"2000";
    tmp(54800) := x"2000";
    tmp(54801) := x"2000";
    tmp(54802) := x"2000";
    tmp(54803) := x"2000";
    tmp(54804) := x"1800";
    tmp(54805) := x"1800";
    tmp(54806) := x"1800";
    tmp(54807) := x"1000";
    tmp(54808) := x"0800";
    tmp(54809) := x"0800";
    tmp(54810) := x"0800";
    tmp(54811) := x"0800";
    tmp(54812) := x"0800";
    tmp(54813) := x"0800";
    tmp(54814) := x"1000";
    tmp(54815) := x"1800";
    tmp(54816) := x"2800";
    tmp(54817) := x"3000";
    tmp(54818) := x"2800";
    tmp(54819) := x"2000";
    tmp(54820) := x"2000";
    tmp(54821) := x"2000";
    tmp(54822) := x"1800";
    tmp(54823) := x"1800";
    tmp(54824) := x"1000";
    tmp(54825) := x"0800";
    tmp(54826) := x"0800";
    tmp(54827) := x"0800";
    tmp(54828) := x"0800";
    tmp(54829) := x"1000";
    tmp(54830) := x"1000";
    tmp(54831) := x"1000";
    tmp(54832) := x"1000";
    tmp(54833) := x"0800";
    tmp(54834) := x"0800";
    tmp(54835) := x"0000";
    tmp(54836) := x"0000";
    tmp(54837) := x"0000";
    tmp(54838) := x"0000";
    tmp(54839) := x"0000";
    tmp(54840) := x"0000";
    tmp(54841) := x"0000";
    tmp(54842) := x"0000";
    tmp(54843) := x"0000";
    tmp(54844) := x"1841";
    tmp(54845) := x"5104";
    tmp(54846) := x"6945";
    tmp(54847) := x"91c8";
    tmp(54848) := x"ba6b";
    tmp(54849) := x"c28d";
    tmp(54850) := x"99ea";
    tmp(54851) := x"8146";
    tmp(54852) := x"c24b";
    tmp(54853) := x"d2ee";
    tmp(54854) := x"9a0a";
    tmp(54855) := x"ba6b";
    tmp(54856) := x"60a3";
    tmp(54857) := x"58a2";
    tmp(54858) := x"c2ec";
    tmp(54859) := x"fd37";
    tmp(54860) := x"99e8";
    tmp(54861) := x"9987";
    tmp(54862) := x"78c4";
    tmp(54863) := x"78e4";
    tmp(54864) := x"daed";
    tmp(54865) := x"b209";
    tmp(54866) := x"3820";
    tmp(54867) := x"5021";
    tmp(54868) := x"7904";
    tmp(54869) := x"f432";
    tmp(54870) := x"3821";
    tmp(54871) := x"8125";
    tmp(54872) := x"f3b0";
    tmp(54873) := x"68a3";
    tmp(54874) := x"7082";
    tmp(54875) := x"7082";
    tmp(54876) := x"9104";
    tmp(54877) := x"3821";
    tmp(54878) := x"3820";
    tmp(54879) := x"70e4";
    tmp(54880) := x"d32d";
    tmp(54881) := x"db4f";
    tmp(54882) := x"ec53";
    tmp(54883) := x"58a2";
    tmp(54884) := x"2000";
    tmp(54885) := x"2800";
    tmp(54886) := x"2800";
    tmp(54887) := x"3000";
    tmp(54888) := x"3800";
    tmp(54889) := x"5800";
    tmp(54890) := x"7800";
    tmp(54891) := x"7000";
    tmp(54892) := x"6800";
    tmp(54893) := x"7800";
    tmp(54894) := x"8800";
    tmp(54895) := x"9020";
    tmp(54896) := x"8000";
    tmp(54897) := x"9020";
    tmp(54898) := x"a820";
    tmp(54899) := x"b020";
    tmp(54900) := x"b820";
    tmp(54901) := x"b820";
    tmp(54902) := x"b820";
    tmp(54903) := x"c020";
    tmp(54904) := x"a800";
    tmp(54905) := x"b820";
    tmp(54906) := x"c020";
    tmp(54907) := x"6840";
    tmp(54908) := x"1020";
    tmp(54909) := x"0820";
    tmp(54910) := x"0840";
    tmp(54911) := x"0840";
    tmp(54912) := x"0820";
    tmp(54913) := x"0840";
    tmp(54914) := x"0820";
    tmp(54915) := x"0820";
    tmp(54916) := x"0820";
    tmp(54917) := x"0820";
    tmp(54918) := x"0820";
    tmp(54919) := x"0840";
    tmp(54920) := x"0840";
    tmp(54921) := x"0840";
    tmp(54922) := x"0840";
    tmp(54923) := x"0840";
    tmp(54924) := x"0840";
    tmp(54925) := x"0840";
    tmp(54926) := x"0840";
    tmp(54927) := x"0840";
    tmp(54928) := x"0840";
    tmp(54929) := x"0840";
    tmp(54930) := x"0840";
    tmp(54931) := x"0840";
    tmp(54932) := x"0840";
    tmp(54933) := x"0840";
    tmp(54934) := x"0820";
    tmp(54935) := x"0820";
    tmp(54936) := x"0820";
    tmp(54937) := x"0820";
    tmp(54938) := x"0820";
    tmp(54939) := x"0820";
    tmp(54940) := x"0820";
    tmp(54941) := x"0820";
    tmp(54942) := x"0820";
    tmp(54943) := x"0820";
    tmp(54944) := x"0820";
    tmp(54945) := x"0820";
    tmp(54946) := x"0820";
    tmp(54947) := x"0820";
    tmp(54948) := x"0820";
    tmp(54949) := x"0820";
    tmp(54950) := x"0820";
    tmp(54951) := x"0820";
    tmp(54952) := x"0820";
    tmp(54953) := x"0820";
    tmp(54954) := x"0820";
    tmp(54955) := x"0820";
    tmp(54956) := x"0820";
    tmp(54957) := x"0820";
    tmp(54958) := x"0820";
    tmp(54959) := x"0820";
    tmp(54960) := x"0000";
    tmp(54961) := x"0000";
    tmp(54962) := x"0000";
    tmp(54963) := x"0800";
    tmp(54964) := x"0800";
    tmp(54965) := x"0800";
    tmp(54966) := x"0800";
    tmp(54967) := x"0800";
    tmp(54968) := x"0800";
    tmp(54969) := x"1000";
    tmp(54970) := x"1000";
    tmp(54971) := x"1000";
    tmp(54972) := x"1000";
    tmp(54973) := x"1000";
    tmp(54974) := x"1800";
    tmp(54975) := x"1800";
    tmp(54976) := x"1000";
    tmp(54977) := x"1800";
    tmp(54978) := x"1800";
    tmp(54979) := x"1800";
    tmp(54980) := x"1800";
    tmp(54981) := x"1800";
    tmp(54982) := x"1800";
    tmp(54983) := x"1800";
    tmp(54984) := x"1800";
    tmp(54985) := x"1800";
    tmp(54986) := x"1800";
    tmp(54987) := x"1800";
    tmp(54988) := x"1800";
    tmp(54989) := x"1800";
    tmp(54990) := x"1800";
    tmp(54991) := x"2000";
    tmp(54992) := x"2000";
    tmp(54993) := x"2000";
    tmp(54994) := x"2000";
    tmp(54995) := x"2000";
    tmp(54996) := x"2000";
    tmp(54997) := x"2000";
    tmp(54998) := x"2000";
    tmp(54999) := x"2800";
    tmp(55000) := x"2800";
    tmp(55001) := x"3000";
    tmp(55002) := x"3000";
    tmp(55003) := x"3000";
    tmp(55004) := x"2800";
    tmp(55005) := x"2800";
    tmp(55006) := x"2800";
    tmp(55007) := x"2800";
    tmp(55008) := x"2800";
    tmp(55009) := x"2800";
    tmp(55010) := x"2800";
    tmp(55011) := x"2800";
    tmp(55012) := x"2800";
    tmp(55013) := x"2800";
    tmp(55014) := x"2800";
    tmp(55015) := x"2800";
    tmp(55016) := x"2800";
    tmp(55017) := x"3000";
    tmp(55018) := x"3000";
    tmp(55019) := x"3000";
    tmp(55020) := x"3800";
    tmp(55021) := x"3800";
    tmp(55022) := x"3800";
    tmp(55023) := x"3000";
    tmp(55024) := x"2800";
    tmp(55025) := x"2800";
    tmp(55026) := x"2800";
    tmp(55027) := x"2000";
    tmp(55028) := x"2000";
    tmp(55029) := x"1800";
    tmp(55030) := x"1800";
    tmp(55031) := x"1000";
    tmp(55032) := x"1000";
    tmp(55033) := x"1000";
    tmp(55034) := x"1800";
    tmp(55035) := x"1800";
    tmp(55036) := x"1800";
    tmp(55037) := x"1800";
    tmp(55038) := x"2000";
    tmp(55039) := x"2000";
    tmp(55040) := x"2800";
    tmp(55041) := x"2000";
    tmp(55042) := x"2000";
    tmp(55043) := x"2000";
    tmp(55044) := x"2000";
    tmp(55045) := x"1800";
    tmp(55046) := x"1800";
    tmp(55047) := x"1800";
    tmp(55048) := x"1000";
    tmp(55049) := x"1000";
    tmp(55050) := x"1000";
    tmp(55051) := x"0800";
    tmp(55052) := x"1000";
    tmp(55053) := x"1000";
    tmp(55054) := x"0800";
    tmp(55055) := x"1000";
    tmp(55056) := x"2800";
    tmp(55057) := x"3800";
    tmp(55058) := x"3820";
    tmp(55059) := x"3820";
    tmp(55060) := x"3000";
    tmp(55061) := x"2800";
    tmp(55062) := x"2000";
    tmp(55063) := x"1800";
    tmp(55064) := x"1000";
    tmp(55065) := x"1000";
    tmp(55066) := x"0800";
    tmp(55067) := x"0800";
    tmp(55068) := x"1000";
    tmp(55069) := x"1800";
    tmp(55070) := x"2000";
    tmp(55071) := x"2800";
    tmp(55072) := x"2800";
    tmp(55073) := x"2000";
    tmp(55074) := x"1800";
    tmp(55075) := x"1000";
    tmp(55076) := x"0800";
    tmp(55077) := x"0000";
    tmp(55078) := x"0000";
    tmp(55079) := x"0000";
    tmp(55080) := x"0000";
    tmp(55081) := x"0000";
    tmp(55082) := x"0000";
    tmp(55083) := x"1861";
    tmp(55084) := x"5104";
    tmp(55085) := x"81c7";
    tmp(55086) := x"99e8";
    tmp(55087) := x"aa2a";
    tmp(55088) := x"b24b";
    tmp(55089) := x"b26c";
    tmp(55090) := x"8187";
    tmp(55091) := x"c24b";
    tmp(55092) := x"ba0a";
    tmp(55093) := x"eaee";
    tmp(55094) := x"b24a";
    tmp(55095) := x"91c8";
    tmp(55096) := x"aa29";
    tmp(55097) := x"6925";
    tmp(55098) := x"9a09";
    tmp(55099) := x"baac";
    tmp(55100) := x"5882";
    tmp(55101) := x"c208";
    tmp(55102) := x"78c4";
    tmp(55103) := x"9166";
    tmp(55104) := x"c22a";
    tmp(55105) := x"a987";
    tmp(55106) := x"4021";
    tmp(55107) := x"6041";
    tmp(55108) := x"4021";
    tmp(55109) := x"e2cc";
    tmp(55110) := x"c24a";
    tmp(55111) := x"3821";
    tmp(55112) := x"8925";
    tmp(55113) := x"c1e8";
    tmp(55114) := x"5021";
    tmp(55115) := x"6841";
    tmp(55116) := x"90c3";
    tmp(55117) := x"88c3";
    tmp(55118) := x"6882";
    tmp(55119) := x"4041";
    tmp(55120) := x"9966";
    tmp(55121) := x"e2ec";
    tmp(55122) := x"f3af";
    tmp(55123) := x"2820";
    tmp(55124) := x"2000";
    tmp(55125) := x"2800";
    tmp(55126) := x"2800";
    tmp(55127) := x"3000";
    tmp(55128) := x"4000";
    tmp(55129) := x"6000";
    tmp(55130) := x"6800";
    tmp(55131) := x"6800";
    tmp(55132) := x"7000";
    tmp(55133) := x"7800";
    tmp(55134) := x"8800";
    tmp(55135) := x"8800";
    tmp(55136) := x"8820";
    tmp(55137) := x"9020";
    tmp(55138) := x"a020";
    tmp(55139) := x"a000";
    tmp(55140) := x"b820";
    tmp(55141) := x"c020";
    tmp(55142) := x"c820";
    tmp(55143) := x"b000";
    tmp(55144) := x"b000";
    tmp(55145) := x"c020";
    tmp(55146) := x"d020";
    tmp(55147) := x"6040";
    tmp(55148) := x"1020";
    tmp(55149) := x"0840";
    tmp(55150) := x"0840";
    tmp(55151) := x"0840";
    tmp(55152) := x"0840";
    tmp(55153) := x"0840";
    tmp(55154) := x"0840";
    tmp(55155) := x"0840";
    tmp(55156) := x"0840";
    tmp(55157) := x"0840";
    tmp(55158) := x"0840";
    tmp(55159) := x"0840";
    tmp(55160) := x"0840";
    tmp(55161) := x"0840";
    tmp(55162) := x"0840";
    tmp(55163) := x"0840";
    tmp(55164) := x"0820";
    tmp(55165) := x"0840";
    tmp(55166) := x"0820";
    tmp(55167) := x"0820";
    tmp(55168) := x"0820";
    tmp(55169) := x"0840";
    tmp(55170) := x"0840";
    tmp(55171) := x"0840";
    tmp(55172) := x"0820";
    tmp(55173) := x"0820";
    tmp(55174) := x"0820";
    tmp(55175) := x"0820";
    tmp(55176) := x"0820";
    tmp(55177) := x"0820";
    tmp(55178) := x"0820";
    tmp(55179) := x"0820";
    tmp(55180) := x"0820";
    tmp(55181) := x"0820";
    tmp(55182) := x"0820";
    tmp(55183) := x"0820";
    tmp(55184) := x"0820";
    tmp(55185) := x"0820";
    tmp(55186) := x"0820";
    tmp(55187) := x"0820";
    tmp(55188) := x"0820";
    tmp(55189) := x"0820";
    tmp(55190) := x"0820";
    tmp(55191) := x"0820";
    tmp(55192) := x"0820";
    tmp(55193) := x"0820";
    tmp(55194) := x"0820";
    tmp(55195) := x"0820";
    tmp(55196) := x"0820";
    tmp(55197) := x"0820";
    tmp(55198) := x"0820";
    tmp(55199) := x"0820";
    tmp(55200) := x"0000";
    tmp(55201) := x"0800";
    tmp(55202) := x"0800";
    tmp(55203) := x"0800";
    tmp(55204) := x"0800";
    tmp(55205) := x"0800";
    tmp(55206) := x"0800";
    tmp(55207) := x"1000";
    tmp(55208) := x"1000";
    tmp(55209) := x"1000";
    tmp(55210) := x"1000";
    tmp(55211) := x"1800";
    tmp(55212) := x"1800";
    tmp(55213) := x"1800";
    tmp(55214) := x"1800";
    tmp(55215) := x"1800";
    tmp(55216) := x"1800";
    tmp(55217) := x"1800";
    tmp(55218) := x"1800";
    tmp(55219) := x"1800";
    tmp(55220) := x"1800";
    tmp(55221) := x"1800";
    tmp(55222) := x"1800";
    tmp(55223) := x"1800";
    tmp(55224) := x"1000";
    tmp(55225) := x"1800";
    tmp(55226) := x"1800";
    tmp(55227) := x"1000";
    tmp(55228) := x"1800";
    tmp(55229) := x"1800";
    tmp(55230) := x"2000";
    tmp(55231) := x"2000";
    tmp(55232) := x"2820";
    tmp(55233) := x"2800";
    tmp(55234) := x"2000";
    tmp(55235) := x"2000";
    tmp(55236) := x"2000";
    tmp(55237) := x"2000";
    tmp(55238) := x"2000";
    tmp(55239) := x"2800";
    tmp(55240) := x"2800";
    tmp(55241) := x"2800";
    tmp(55242) := x"3000";
    tmp(55243) := x"2800";
    tmp(55244) := x"2800";
    tmp(55245) := x"2800";
    tmp(55246) := x"2800";
    tmp(55247) := x"2000";
    tmp(55248) := x"2800";
    tmp(55249) := x"2800";
    tmp(55250) := x"2800";
    tmp(55251) := x"2800";
    tmp(55252) := x"2800";
    tmp(55253) := x"2800";
    tmp(55254) := x"2800";
    tmp(55255) := x"2800";
    tmp(55256) := x"2800";
    tmp(55257) := x"3000";
    tmp(55258) := x"3000";
    tmp(55259) := x"3800";
    tmp(55260) := x"3800";
    tmp(55261) := x"3800";
    tmp(55262) := x"3800";
    tmp(55263) := x"3000";
    tmp(55264) := x"2800";
    tmp(55265) := x"2800";
    tmp(55266) := x"2800";
    tmp(55267) := x"2000";
    tmp(55268) := x"2000";
    tmp(55269) := x"2000";
    tmp(55270) := x"2000";
    tmp(55271) := x"1800";
    tmp(55272) := x"1000";
    tmp(55273) := x"1000";
    tmp(55274) := x"1800";
    tmp(55275) := x"1800";
    tmp(55276) := x"1800";
    tmp(55277) := x"2000";
    tmp(55278) := x"2000";
    tmp(55279) := x"2800";
    tmp(55280) := x"2800";
    tmp(55281) := x"2800";
    tmp(55282) := x"2800";
    tmp(55283) := x"2800";
    tmp(55284) := x"2000";
    tmp(55285) := x"2000";
    tmp(55286) := x"1800";
    tmp(55287) := x"1000";
    tmp(55288) := x"1800";
    tmp(55289) := x"1800";
    tmp(55290) := x"1800";
    tmp(55291) := x"1800";
    tmp(55292) := x"1800";
    tmp(55293) := x"1000";
    tmp(55294) := x"1000";
    tmp(55295) := x"0800";
    tmp(55296) := x"1000";
    tmp(55297) := x"1000";
    tmp(55298) := x"1800";
    tmp(55299) := x"2000";
    tmp(55300) := x"2000";
    tmp(55301) := x"2000";
    tmp(55302) := x"2800";
    tmp(55303) := x"2800";
    tmp(55304) := x"2800";
    tmp(55305) := x"2800";
    tmp(55306) := x"2020";
    tmp(55307) := x"1800";
    tmp(55308) := x"2000";
    tmp(55309) := x"2000";
    tmp(55310) := x"2800";
    tmp(55311) := x"3000";
    tmp(55312) := x"3020";
    tmp(55313) := x"3020";
    tmp(55314) := x"3020";
    tmp(55315) := x"2820";
    tmp(55316) := x"2020";
    tmp(55317) := x"0800";
    tmp(55318) := x"0000";
    tmp(55319) := x"0000";
    tmp(55320) := x"0000";
    tmp(55321) := x"0000";
    tmp(55322) := x"2061";
    tmp(55323) := x"5104";
    tmp(55324) := x"89c7";
    tmp(55325) := x"aa6a";
    tmp(55326) := x"99e9";
    tmp(55327) := x"99e9";
    tmp(55328) := x"9a0a";
    tmp(55329) := x"99e9";
    tmp(55330) := x"6905";
    tmp(55331) := x"b20a";
    tmp(55332) := x"b1ea";
    tmp(55333) := x"a1a8";
    tmp(55334) := x"8987";
    tmp(55335) := x"a209";
    tmp(55336) := x"db4f";
    tmp(55337) := x"7166";
    tmp(55338) := x"db2d";
    tmp(55339) := x"a1a7";
    tmp(55340) := x"5041";
    tmp(55341) := x"fb6e";
    tmp(55342) := x"78e4";
    tmp(55343) := x"9125";
    tmp(55344) := x"9925";
    tmp(55345) := x"9146";
    tmp(55346) := x"70a3";
    tmp(55347) := x"7061";
    tmp(55348) := x"3000";
    tmp(55349) := x"70a2";
    tmp(55350) := x"f3ae";
    tmp(55351) := x"aa4a";
    tmp(55352) := x"4020";
    tmp(55353) := x"a104";
    tmp(55354) := x"a0e3";
    tmp(55355) := x"5821";
    tmp(55356) := x"6841";
    tmp(55357) := x"7062";
    tmp(55358) := x"6061";
    tmp(55359) := x"78a2";
    tmp(55360) := x"5041";
    tmp(55361) := x"78c3";
    tmp(55362) := x"b9c6";
    tmp(55363) := x"2000";
    tmp(55364) := x"2800";
    tmp(55365) := x"3000";
    tmp(55366) := x"2800";
    tmp(55367) := x"3000";
    tmp(55368) := x"4800";
    tmp(55369) := x"6800";
    tmp(55370) := x"7000";
    tmp(55371) := x"7000";
    tmp(55372) := x"8000";
    tmp(55373) := x"8800";
    tmp(55374) := x"8800";
    tmp(55375) := x"9000";
    tmp(55376) := x"9820";
    tmp(55377) := x"a020";
    tmp(55378) := x"a820";
    tmp(55379) := x"a000";
    tmp(55380) := x"c820";
    tmp(55381) := x"b820";
    tmp(55382) := x"b820";
    tmp(55383) := x"b000";
    tmp(55384) := x"b000";
    tmp(55385) := x"d820";
    tmp(55386) := x"d840";
    tmp(55387) := x"5840";
    tmp(55388) := x"1040";
    tmp(55389) := x"0840";
    tmp(55390) := x"0840";
    tmp(55391) := x"0840";
    tmp(55392) := x"0840";
    tmp(55393) := x"0840";
    tmp(55394) := x"0840";
    tmp(55395) := x"0840";
    tmp(55396) := x"0840";
    tmp(55397) := x"0840";
    tmp(55398) := x"0840";
    tmp(55399) := x"0840";
    tmp(55400) := x"0840";
    tmp(55401) := x"0840";
    tmp(55402) := x"0840";
    tmp(55403) := x"0840";
    tmp(55404) := x"0840";
    tmp(55405) := x"0820";
    tmp(55406) := x"0820";
    tmp(55407) := x"0840";
    tmp(55408) := x"0840";
    tmp(55409) := x"0840";
    tmp(55410) := x"0820";
    tmp(55411) := x"0820";
    tmp(55412) := x"0820";
    tmp(55413) := x"0820";
    tmp(55414) := x"0820";
    tmp(55415) := x"0820";
    tmp(55416) := x"0820";
    tmp(55417) := x"0820";
    tmp(55418) := x"0820";
    tmp(55419) := x"0820";
    tmp(55420) := x"0820";
    tmp(55421) := x"0820";
    tmp(55422) := x"0820";
    tmp(55423) := x"0820";
    tmp(55424) := x"0820";
    tmp(55425) := x"0820";
    tmp(55426) := x"0820";
    tmp(55427) := x"0820";
    tmp(55428) := x"0820";
    tmp(55429) := x"0820";
    tmp(55430) := x"0820";
    tmp(55431) := x"0820";
    tmp(55432) := x"0820";
    tmp(55433) := x"0820";
    tmp(55434) := x"0820";
    tmp(55435) := x"0820";
    tmp(55436) := x"0820";
    tmp(55437) := x"0820";
    tmp(55438) := x"0820";
    tmp(55439) := x"0820";
    tmp(55440) := x"0000";
    tmp(55441) := x"0800";
    tmp(55442) := x"0800";
    tmp(55443) := x"0800";
    tmp(55444) := x"0800";
    tmp(55445) := x"1000";
    tmp(55446) := x"1000";
    tmp(55447) := x"1000";
    tmp(55448) := x"1000";
    tmp(55449) := x"1000";
    tmp(55450) := x"1000";
    tmp(55451) := x"1000";
    tmp(55452) := x"1800";
    tmp(55453) := x"1800";
    tmp(55454) := x"1800";
    tmp(55455) := x"1800";
    tmp(55456) := x"1800";
    tmp(55457) := x"1000";
    tmp(55458) := x"1000";
    tmp(55459) := x"1000";
    tmp(55460) := x"1800";
    tmp(55461) := x"1800";
    tmp(55462) := x"1800";
    tmp(55463) := x"1800";
    tmp(55464) := x"1800";
    tmp(55465) := x"1800";
    tmp(55466) := x"1800";
    tmp(55467) := x"1800";
    tmp(55468) := x"2000";
    tmp(55469) := x"2000";
    tmp(55470) := x"2000";
    tmp(55471) := x"2800";
    tmp(55472) := x"2800";
    tmp(55473) := x"2000";
    tmp(55474) := x"2000";
    tmp(55475) := x"2000";
    tmp(55476) := x"2000";
    tmp(55477) := x"2000";
    tmp(55478) := x"2000";
    tmp(55479) := x"2000";
    tmp(55480) := x"2000";
    tmp(55481) := x"2800";
    tmp(55482) := x"2800";
    tmp(55483) := x"2800";
    tmp(55484) := x"2800";
    tmp(55485) := x"2800";
    tmp(55486) := x"2800";
    tmp(55487) := x"2800";
    tmp(55488) := x"2800";
    tmp(55489) := x"2800";
    tmp(55490) := x"2800";
    tmp(55491) := x"2800";
    tmp(55492) := x"2800";
    tmp(55493) := x"2800";
    tmp(55494) := x"3000";
    tmp(55495) := x"3000";
    tmp(55496) := x"2800";
    tmp(55497) := x"2800";
    tmp(55498) := x"3000";
    tmp(55499) := x"3000";
    tmp(55500) := x"3800";
    tmp(55501) := x"3800";
    tmp(55502) := x"3800";
    tmp(55503) := x"3800";
    tmp(55504) := x"3000";
    tmp(55505) := x"2800";
    tmp(55506) := x"2800";
    tmp(55507) := x"2000";
    tmp(55508) := x"2800";
    tmp(55509) := x"2800";
    tmp(55510) := x"2000";
    tmp(55511) := x"2000";
    tmp(55512) := x"1800";
    tmp(55513) := x"1000";
    tmp(55514) := x"1000";
    tmp(55515) := x"1800";
    tmp(55516) := x"1800";
    tmp(55517) := x"2000";
    tmp(55518) := x"2000";
    tmp(55519) := x"2800";
    tmp(55520) := x"2800";
    tmp(55521) := x"2800";
    tmp(55522) := x"2800";
    tmp(55523) := x"2800";
    tmp(55524) := x"2820";
    tmp(55525) := x"2820";
    tmp(55526) := x"1800";
    tmp(55527) := x"1800";
    tmp(55528) := x"1800";
    tmp(55529) := x"1800";
    tmp(55530) := x"2000";
    tmp(55531) := x"2000";
    tmp(55532) := x"2000";
    tmp(55533) := x"1800";
    tmp(55534) := x"1000";
    tmp(55535) := x"1000";
    tmp(55536) := x"0800";
    tmp(55537) := x"0800";
    tmp(55538) := x"0800";
    tmp(55539) := x"1000";
    tmp(55540) := x"1800";
    tmp(55541) := x"2000";
    tmp(55542) := x"2800";
    tmp(55543) := x"3000";
    tmp(55544) := x"2800";
    tmp(55545) := x"2800";
    tmp(55546) := x"3000";
    tmp(55547) := x"2800";
    tmp(55548) := x"2800";
    tmp(55549) := x"3000";
    tmp(55550) := x"3800";
    tmp(55551) := x"3800";
    tmp(55552) := x"3820";
    tmp(55553) := x"3020";
    tmp(55554) := x"3020";
    tmp(55555) := x"3020";
    tmp(55556) := x"3020";
    tmp(55557) := x"2820";
    tmp(55558) := x"1020";
    tmp(55559) := x"0000";
    tmp(55560) := x"0820";
    tmp(55561) := x"28a2";
    tmp(55562) := x"48e3";
    tmp(55563) := x"79c7";
    tmp(55564) := x"6145";
    tmp(55565) := x"6925";
    tmp(55566) := x"8187";
    tmp(55567) := x"7946";
    tmp(55568) := x"7966";
    tmp(55569) := x"6925";
    tmp(55570) := x"8166";
    tmp(55571) := x"c26b";
    tmp(55572) := x"ba2a";
    tmp(55573) := x"b20a";
    tmp(55574) := x"d2ad";
    tmp(55575) := x"89a8";
    tmp(55576) := x"b26b";
    tmp(55577) := x"7145";
    tmp(55578) := x"ebf0";
    tmp(55579) := x"b209";
    tmp(55580) := x"5861";
    tmp(55581) := x"f3cf";
    tmp(55582) := x"68e4";
    tmp(55583) := x"78c4";
    tmp(55584) := x"80c3";
    tmp(55585) := x"70a3";
    tmp(55586) := x"a1a8";
    tmp(55587) := x"4021";
    tmp(55588) := x"4820";
    tmp(55589) := x"4820";
    tmp(55590) := x"70a3";
    tmp(55591) := x"dbaf";
    tmp(55592) := x"7882";
    tmp(55593) := x"5841";
    tmp(55594) := x"eacb";
    tmp(55595) := x"7061";
    tmp(55596) := x"7861";
    tmp(55597) := x"6041";
    tmp(55598) := x"4000";
    tmp(55599) := x"6041";
    tmp(55600) := x"6861";
    tmp(55601) := x"5041";
    tmp(55602) := x"6061";
    tmp(55603) := x"2000";
    tmp(55604) := x"2800";
    tmp(55605) := x"2800";
    tmp(55606) := x"2800";
    tmp(55607) := x"3800";
    tmp(55608) := x"5800";
    tmp(55609) := x"7000";
    tmp(55610) := x"6800";
    tmp(55611) := x"7000";
    tmp(55612) := x"8800";
    tmp(55613) := x"8820";
    tmp(55614) := x"7800";
    tmp(55615) := x"8800";
    tmp(55616) := x"9820";
    tmp(55617) := x"9820";
    tmp(55618) := x"9800";
    tmp(55619) := x"9800";
    tmp(55620) := x"a000";
    tmp(55621) := x"b000";
    tmp(55622) := x"b000";
    tmp(55623) := x"b000";
    tmp(55624) := x"b000";
    tmp(55625) := x"d820";
    tmp(55626) := x"c840";
    tmp(55627) := x"4040";
    tmp(55628) := x"1040";
    tmp(55629) := x"0841";
    tmp(55630) := x"0841";
    tmp(55631) := x"0840";
    tmp(55632) := x"0840";
    tmp(55633) := x"0841";
    tmp(55634) := x"0840";
    tmp(55635) := x"0840";
    tmp(55636) := x"0840";
    tmp(55637) := x"0840";
    tmp(55638) := x"0840";
    tmp(55639) := x"0840";
    tmp(55640) := x"0840";
    tmp(55641) := x"0840";
    tmp(55642) := x"0840";
    tmp(55643) := x"0840";
    tmp(55644) := x"0840";
    tmp(55645) := x"0820";
    tmp(55646) := x"0820";
    tmp(55647) := x"0820";
    tmp(55648) := x"0820";
    tmp(55649) := x"0840";
    tmp(55650) := x"0820";
    tmp(55651) := x"0820";
    tmp(55652) := x"0820";
    tmp(55653) := x"0820";
    tmp(55654) := x"0820";
    tmp(55655) := x"0820";
    tmp(55656) := x"0820";
    tmp(55657) := x"0820";
    tmp(55658) := x"0820";
    tmp(55659) := x"0820";
    tmp(55660) := x"0820";
    tmp(55661) := x"0820";
    tmp(55662) := x"0820";
    tmp(55663) := x"0820";
    tmp(55664) := x"0820";
    tmp(55665) := x"0820";
    tmp(55666) := x"0820";
    tmp(55667) := x"0820";
    tmp(55668) := x"0820";
    tmp(55669) := x"0820";
    tmp(55670) := x"0820";
    tmp(55671) := x"0820";
    tmp(55672) := x"0820";
    tmp(55673) := x"0820";
    tmp(55674) := x"0820";
    tmp(55675) := x"0820";
    tmp(55676) := x"0820";
    tmp(55677) := x"0820";
    tmp(55678) := x"0820";
    tmp(55679) := x"0820";
    tmp(55680) := x"0000";
    tmp(55681) := x"0800";
    tmp(55682) := x"0800";
    tmp(55683) := x"0800";
    tmp(55684) := x"1000";
    tmp(55685) := x"1000";
    tmp(55686) := x"1000";
    tmp(55687) := x"1000";
    tmp(55688) := x"1000";
    tmp(55689) := x"1000";
    tmp(55690) := x"1800";
    tmp(55691) := x"1800";
    tmp(55692) := x"1800";
    tmp(55693) := x"1800";
    tmp(55694) := x"1000";
    tmp(55695) := x"1000";
    tmp(55696) := x"1000";
    tmp(55697) := x"1000";
    tmp(55698) := x"1000";
    tmp(55699) := x"1800";
    tmp(55700) := x"1800";
    tmp(55701) := x"1800";
    tmp(55702) := x"1800";
    tmp(55703) := x"1800";
    tmp(55704) := x"1800";
    tmp(55705) := x"2000";
    tmp(55706) := x"2000";
    tmp(55707) := x"2000";
    tmp(55708) := x"2000";
    tmp(55709) := x"2000";
    tmp(55710) := x"2000";
    tmp(55711) := x"2800";
    tmp(55712) := x"2800";
    tmp(55713) := x"2800";
    tmp(55714) := x"2000";
    tmp(55715) := x"2000";
    tmp(55716) := x"2000";
    tmp(55717) := x"2000";
    tmp(55718) := x"2000";
    tmp(55719) := x"2800";
    tmp(55720) := x"2000";
    tmp(55721) := x"2800";
    tmp(55722) := x"2800";
    tmp(55723) := x"3000";
    tmp(55724) := x"2800";
    tmp(55725) := x"2800";
    tmp(55726) := x"2800";
    tmp(55727) := x"2800";
    tmp(55728) := x"2800";
    tmp(55729) := x"2800";
    tmp(55730) := x"2800";
    tmp(55731) := x"2800";
    tmp(55732) := x"2800";
    tmp(55733) := x"2800";
    tmp(55734) := x"3000";
    tmp(55735) := x"3000";
    tmp(55736) := x"3000";
    tmp(55737) := x"3000";
    tmp(55738) := x"2800";
    tmp(55739) := x"3000";
    tmp(55740) := x"3000";
    tmp(55741) := x"3000";
    tmp(55742) := x"2800";
    tmp(55743) := x"2000";
    tmp(55744) := x"1800";
    tmp(55745) := x"1800";
    tmp(55746) := x"2000";
    tmp(55747) := x"2000";
    tmp(55748) := x"2000";
    tmp(55749) := x"2800";
    tmp(55750) := x"2000";
    tmp(55751) := x"2000";
    tmp(55752) := x"2000";
    tmp(55753) := x"1800";
    tmp(55754) := x"1800";
    tmp(55755) := x"1800";
    tmp(55756) := x"1800";
    tmp(55757) := x"1800";
    tmp(55758) := x"2000";
    tmp(55759) := x"2000";
    tmp(55760) := x"2800";
    tmp(55761) := x"2800";
    tmp(55762) := x"2800";
    tmp(55763) := x"3020";
    tmp(55764) := x"3020";
    tmp(55765) := x"2820";
    tmp(55766) := x"2000";
    tmp(55767) := x"1800";
    tmp(55768) := x"1800";
    tmp(55769) := x"2000";
    tmp(55770) := x"2000";
    tmp(55771) := x"2800";
    tmp(55772) := x"2000";
    tmp(55773) := x"1800";
    tmp(55774) := x"1800";
    tmp(55775) := x"1000";
    tmp(55776) := x"0800";
    tmp(55777) := x"0800";
    tmp(55778) := x"1000";
    tmp(55779) := x"1800";
    tmp(55780) := x"2000";
    tmp(55781) := x"2000";
    tmp(55782) := x"2800";
    tmp(55783) := x"3000";
    tmp(55784) := x"2800";
    tmp(55785) := x"3000";
    tmp(55786) := x"3000";
    tmp(55787) := x"3000";
    tmp(55788) := x"3800";
    tmp(55789) := x"3800";
    tmp(55790) := x"4000";
    tmp(55791) := x"4800";
    tmp(55792) := x"4820";
    tmp(55793) := x"4020";
    tmp(55794) := x"4020";
    tmp(55795) := x"3820";
    tmp(55796) := x"3020";
    tmp(55797) := x"2820";
    tmp(55798) := x"2020";
    tmp(55799) := x"1020";
    tmp(55800) := x"1841";
    tmp(55801) := x"30a2";
    tmp(55802) := x"40c3";
    tmp(55803) := x"48e4";
    tmp(55804) := x"48c4";
    tmp(55805) := x"7146";
    tmp(55806) := x"8166";
    tmp(55807) := x"8146";
    tmp(55808) := x"8166";
    tmp(55809) := x"7125";
    tmp(55810) := x"8966";
    tmp(55811) := x"8967";
    tmp(55812) := x"ca8c";
    tmp(55813) := x"99c8";
    tmp(55814) := x"b24a";
    tmp(55815) := x"a1e9";
    tmp(55816) := x"b1c8";
    tmp(55817) := x"4041";
    tmp(55818) := x"c24a";
    tmp(55819) := x"9125";
    tmp(55820) := x"5041";
    tmp(55821) := x"eacb";
    tmp(55822) := x"78c4";
    tmp(55823) := x"9966";
    tmp(55824) := x"78c3";
    tmp(55825) := x"6061";
    tmp(55826) := x"ebb0";
    tmp(55827) := x"4041";
    tmp(55828) := x"6041";
    tmp(55829) := x"6821";
    tmp(55830) := x"6841";
    tmp(55831) := x"9125";
    tmp(55832) := x"da08";
    tmp(55833) := x"5821";
    tmp(55834) := x"b166";
    tmp(55835) := x"8882";
    tmp(55836) := x"a0e4";
    tmp(55837) := x"88a3";
    tmp(55838) := x"5020";
    tmp(55839) := x"5020";
    tmp(55840) := x"88a2";
    tmp(55841) := x"5841";
    tmp(55842) := x"3020";
    tmp(55843) := x"2800";
    tmp(55844) := x"3000";
    tmp(55845) := x"2000";
    tmp(55846) := x"2800";
    tmp(55847) := x"4800";
    tmp(55848) := x"6000";
    tmp(55849) := x"6000";
    tmp(55850) := x"6000";
    tmp(55851) := x"7000";
    tmp(55852) := x"8800";
    tmp(55853) := x"8800";
    tmp(55854) := x"8800";
    tmp(55855) := x"8000";
    tmp(55856) := x"9800";
    tmp(55857) := x"9000";
    tmp(55858) := x"9000";
    tmp(55859) := x"9000";
    tmp(55860) := x"9800";
    tmp(55861) := x"a800";
    tmp(55862) := x"b820";
    tmp(55863) := x"b000";
    tmp(55864) := x"b820";
    tmp(55865) := x"c820";
    tmp(55866) := x"b840";
    tmp(55867) := x"3040";
    tmp(55868) := x"0840";
    tmp(55869) := x"0841";
    tmp(55870) := x"0841";
    tmp(55871) := x"0840";
    tmp(55872) := x"0841";
    tmp(55873) := x"0841";
    tmp(55874) := x"0840";
    tmp(55875) := x"0840";
    tmp(55876) := x"0840";
    tmp(55877) := x"0840";
    tmp(55878) := x"0840";
    tmp(55879) := x"0840";
    tmp(55880) := x"0840";
    tmp(55881) := x"0840";
    tmp(55882) := x"0840";
    tmp(55883) := x"0840";
    tmp(55884) := x"0840";
    tmp(55885) := x"0820";
    tmp(55886) := x"0820";
    tmp(55887) := x"0820";
    tmp(55888) := x"0820";
    tmp(55889) := x"0820";
    tmp(55890) := x"0820";
    tmp(55891) := x"0820";
    tmp(55892) := x"0820";
    tmp(55893) := x"0820";
    tmp(55894) := x"0820";
    tmp(55895) := x"0820";
    tmp(55896) := x"0820";
    tmp(55897) := x"0820";
    tmp(55898) := x"0820";
    tmp(55899) := x"0820";
    tmp(55900) := x"0820";
    tmp(55901) := x"0820";
    tmp(55902) := x"0820";
    tmp(55903) := x"0820";
    tmp(55904) := x"0820";
    tmp(55905) := x"0820";
    tmp(55906) := x"0820";
    tmp(55907) := x"0820";
    tmp(55908) := x"0820";
    tmp(55909) := x"0820";
    tmp(55910) := x"0820";
    tmp(55911) := x"0820";
    tmp(55912) := x"0820";
    tmp(55913) := x"0820";
    tmp(55914) := x"0820";
    tmp(55915) := x"0820";
    tmp(55916) := x"0820";
    tmp(55917) := x"0820";
    tmp(55918) := x"0820";
    tmp(55919) := x"0820";
    tmp(55920) := x"0000";
    tmp(55921) := x"1000";
    tmp(55922) := x"0800";
    tmp(55923) := x"1000";
    tmp(55924) := x"1000";
    tmp(55925) := x"1000";
    tmp(55926) := x"1000";
    tmp(55927) := x"1000";
    tmp(55928) := x"1800";
    tmp(55929) := x"1800";
    tmp(55930) := x"1800";
    tmp(55931) := x"1800";
    tmp(55932) := x"1000";
    tmp(55933) := x"1000";
    tmp(55934) := x"1000";
    tmp(55935) := x"1000";
    tmp(55936) := x"1000";
    tmp(55937) := x"1000";
    tmp(55938) := x"1800";
    tmp(55939) := x"1800";
    tmp(55940) := x"1800";
    tmp(55941) := x"1800";
    tmp(55942) := x"1800";
    tmp(55943) := x"1800";
    tmp(55944) := x"2000";
    tmp(55945) := x"2000";
    tmp(55946) := x"2000";
    tmp(55947) := x"2000";
    tmp(55948) := x"2000";
    tmp(55949) := x"2800";
    tmp(55950) := x"2820";
    tmp(55951) := x"2800";
    tmp(55952) := x"2800";
    tmp(55953) := x"2000";
    tmp(55954) := x"2000";
    tmp(55955) := x"2000";
    tmp(55956) := x"2000";
    tmp(55957) := x"2800";
    tmp(55958) := x"2800";
    tmp(55959) := x"2800";
    tmp(55960) := x"2800";
    tmp(55961) := x"2800";
    tmp(55962) := x"2800";
    tmp(55963) := x"2800";
    tmp(55964) := x"2800";
    tmp(55965) := x"3000";
    tmp(55966) := x"2800";
    tmp(55967) := x"2800";
    tmp(55968) := x"2800";
    tmp(55969) := x"2800";
    tmp(55970) := x"2800";
    tmp(55971) := x"2800";
    tmp(55972) := x"2800";
    tmp(55973) := x"2800";
    tmp(55974) := x"2800";
    tmp(55975) := x"3000";
    tmp(55976) := x"3000";
    tmp(55977) := x"3000";
    tmp(55978) := x"3000";
    tmp(55979) := x"3000";
    tmp(55980) := x"3000";
    tmp(55981) := x"3000";
    tmp(55982) := x"2800";
    tmp(55983) := x"2800";
    tmp(55984) := x"2000";
    tmp(55985) := x"2000";
    tmp(55986) := x"2000";
    tmp(55987) := x"2000";
    tmp(55988) := x"2000";
    tmp(55989) := x"2000";
    tmp(55990) := x"2000";
    tmp(55991) := x"2000";
    tmp(55992) := x"1800";
    tmp(55993) := x"1800";
    tmp(55994) := x"1000";
    tmp(55995) := x"1000";
    tmp(55996) := x"1000";
    tmp(55997) := x"1800";
    tmp(55998) := x"2000";
    tmp(55999) := x"2800";
    tmp(56000) := x"2800";
    tmp(56001) := x"2000";
    tmp(56002) := x"2800";
    tmp(56003) := x"2800";
    tmp(56004) := x"2820";
    tmp(56005) := x"2820";
    tmp(56006) := x"2000";
    tmp(56007) := x"2000";
    tmp(56008) := x"1800";
    tmp(56009) := x"1800";
    tmp(56010) := x"2000";
    tmp(56011) := x"2000";
    tmp(56012) := x"1800";
    tmp(56013) := x"2000";
    tmp(56014) := x"1800";
    tmp(56015) := x"2000";
    tmp(56016) := x"1800";
    tmp(56017) := x"1000";
    tmp(56018) := x"1800";
    tmp(56019) := x"1800";
    tmp(56020) := x"2000";
    tmp(56021) := x"2000";
    tmp(56022) := x"2800";
    tmp(56023) := x"2800";
    tmp(56024) := x"2800";
    tmp(56025) := x"2800";
    tmp(56026) := x"3000";
    tmp(56027) := x"4000";
    tmp(56028) := x"4000";
    tmp(56029) := x"3800";
    tmp(56030) := x"3800";
    tmp(56031) := x"3800";
    tmp(56032) := x"3800";
    tmp(56033) := x"3800";
    tmp(56034) := x"3000";
    tmp(56035) := x"3000";
    tmp(56036) := x"2800";
    tmp(56037) := x"2000";
    tmp(56038) := x"2000";
    tmp(56039) := x"1800";
    tmp(56040) := x"1000";
    tmp(56041) := x"2020";
    tmp(56042) := x"2841";
    tmp(56043) := x"3082";
    tmp(56044) := x"6925";
    tmp(56045) := x"7125";
    tmp(56046) := x"60e4";
    tmp(56047) := x"60e4";
    tmp(56048) := x"6904";
    tmp(56049) := x"58c4";
    tmp(56050) := x"99a8";
    tmp(56051) := x"b24a";
    tmp(56052) := x"8987";
    tmp(56053) := x"b22a";
    tmp(56054) := x"ba6b";
    tmp(56055) := x"91c8";
    tmp(56056) := x"68a2";
    tmp(56057) := x"4841";
    tmp(56058) := x"c1e8";
    tmp(56059) := x"6862";
    tmp(56060) := x"5841";
    tmp(56061) := x"f28a";
    tmp(56062) := x"a166";
    tmp(56063) := x"d24a";
    tmp(56064) := x"6082";
    tmp(56065) := x"6861";
    tmp(56066) := x"ca49";
    tmp(56067) := x"9925";
    tmp(56068) := x"3820";
    tmp(56069) := x"9061";
    tmp(56070) := x"8862";
    tmp(56071) := x"c1e9";
    tmp(56072) := x"80a3";
    tmp(56073) := x"8082";
    tmp(56074) := x"a925";
    tmp(56075) := x"7862";
    tmp(56076) := x"80a2";
    tmp(56077) := x"ea6a";
    tmp(56078) := x"7861";
    tmp(56079) := x"5020";
    tmp(56080) := x"8082";
    tmp(56081) := x"9103";
    tmp(56082) := x"3020";
    tmp(56083) := x"2800";
    tmp(56084) := x"2800";
    tmp(56085) := x"2000";
    tmp(56086) := x"3000";
    tmp(56087) := x"4800";
    tmp(56088) := x"5800";
    tmp(56089) := x"6000";
    tmp(56090) := x"6000";
    tmp(56091) := x"7000";
    tmp(56092) := x"8800";
    tmp(56093) := x"8000";
    tmp(56094) := x"8000";
    tmp(56095) := x"8000";
    tmp(56096) := x"9000";
    tmp(56097) := x"9000";
    tmp(56098) := x"9000";
    tmp(56099) := x"9000";
    tmp(56100) := x"a000";
    tmp(56101) := x"a820";
    tmp(56102) := x"b820";
    tmp(56103) := x"c020";
    tmp(56104) := x"b020";
    tmp(56105) := x"b820";
    tmp(56106) := x"a040";
    tmp(56107) := x"2840";
    tmp(56108) := x"0840";
    tmp(56109) := x"0841";
    tmp(56110) := x"0841";
    tmp(56111) := x"0841";
    tmp(56112) := x"0840";
    tmp(56113) := x"0841";
    tmp(56114) := x"0840";
    tmp(56115) := x"0840";
    tmp(56116) := x"0840";
    tmp(56117) := x"0840";
    tmp(56118) := x"0840";
    tmp(56119) := x"0840";
    tmp(56120) := x"0840";
    tmp(56121) := x"0840";
    tmp(56122) := x"0840";
    tmp(56123) := x"0820";
    tmp(56124) := x"0820";
    tmp(56125) := x"0820";
    tmp(56126) := x"0820";
    tmp(56127) := x"0820";
    tmp(56128) := x"0820";
    tmp(56129) := x"0820";
    tmp(56130) := x"0820";
    tmp(56131) := x"0820";
    tmp(56132) := x"0820";
    tmp(56133) := x"0820";
    tmp(56134) := x"0820";
    tmp(56135) := x"0820";
    tmp(56136) := x"0820";
    tmp(56137) := x"0820";
    tmp(56138) := x"0820";
    tmp(56139) := x"0820";
    tmp(56140) := x"0820";
    tmp(56141) := x"0820";
    tmp(56142) := x"0820";
    tmp(56143) := x"0820";
    tmp(56144) := x"0820";
    tmp(56145) := x"0820";
    tmp(56146) := x"0820";
    tmp(56147) := x"0820";
    tmp(56148) := x"0820";
    tmp(56149) := x"0820";
    tmp(56150) := x"0820";
    tmp(56151) := x"0820";
    tmp(56152) := x"0820";
    tmp(56153) := x"0820";
    tmp(56154) := x"0820";
    tmp(56155) := x"0820";
    tmp(56156) := x"0820";
    tmp(56157) := x"0820";
    tmp(56158) := x"0820";
    tmp(56159) := x"0820";
    tmp(56160) := x"0000";
    tmp(56161) := x"0800";
    tmp(56162) := x"0800";
    tmp(56163) := x"1000";
    tmp(56164) := x"1000";
    tmp(56165) := x"1000";
    tmp(56166) := x"1800";
    tmp(56167) := x"1800";
    tmp(56168) := x"1800";
    tmp(56169) := x"1800";
    tmp(56170) := x"1000";
    tmp(56171) := x"1000";
    tmp(56172) := x"1000";
    tmp(56173) := x"1000";
    tmp(56174) := x"1000";
    tmp(56175) := x"1000";
    tmp(56176) := x"1800";
    tmp(56177) := x"1800";
    tmp(56178) := x"1800";
    tmp(56179) := x"1800";
    tmp(56180) := x"1800";
    tmp(56181) := x"1800";
    tmp(56182) := x"1800";
    tmp(56183) := x"2000";
    tmp(56184) := x"2020";
    tmp(56185) := x"2000";
    tmp(56186) := x"2000";
    tmp(56187) := x"2820";
    tmp(56188) := x"2800";
    tmp(56189) := x"2000";
    tmp(56190) := x"2000";
    tmp(56191) := x"2000";
    tmp(56192) := x"1800";
    tmp(56193) := x"2000";
    tmp(56194) := x"2000";
    tmp(56195) := x"2000";
    tmp(56196) := x"2800";
    tmp(56197) := x"2800";
    tmp(56198) := x"2800";
    tmp(56199) := x"3020";
    tmp(56200) := x"2800";
    tmp(56201) := x"2800";
    tmp(56202) := x"2800";
    tmp(56203) := x"2800";
    tmp(56204) := x"2800";
    tmp(56205) := x"3000";
    tmp(56206) := x"2800";
    tmp(56207) := x"2800";
    tmp(56208) := x"2800";
    tmp(56209) := x"3000";
    tmp(56210) := x"2800";
    tmp(56211) := x"2800";
    tmp(56212) := x"2800";
    tmp(56213) := x"2800";
    tmp(56214) := x"3000";
    tmp(56215) := x"2800";
    tmp(56216) := x"3000";
    tmp(56217) := x"3000";
    tmp(56218) := x"3000";
    tmp(56219) := x"3000";
    tmp(56220) := x"3000";
    tmp(56221) := x"3800";
    tmp(56222) := x"3800";
    tmp(56223) := x"3000";
    tmp(56224) := x"2800";
    tmp(56225) := x"2800";
    tmp(56226) := x"2800";
    tmp(56227) := x"2000";
    tmp(56228) := x"2000";
    tmp(56229) := x"2800";
    tmp(56230) := x"2000";
    tmp(56231) := x"2000";
    tmp(56232) := x"1800";
    tmp(56233) := x"1800";
    tmp(56234) := x"1000";
    tmp(56235) := x"1000";
    tmp(56236) := x"1000";
    tmp(56237) := x"1800";
    tmp(56238) := x"2000";
    tmp(56239) := x"2000";
    tmp(56240) := x"2800";
    tmp(56241) := x"2800";
    tmp(56242) := x"2800";
    tmp(56243) := x"2000";
    tmp(56244) := x"2800";
    tmp(56245) := x"2000";
    tmp(56246) := x"2000";
    tmp(56247) := x"2000";
    tmp(56248) := x"1800";
    tmp(56249) := x"1000";
    tmp(56250) := x"1800";
    tmp(56251) := x"1800";
    tmp(56252) := x"2000";
    tmp(56253) := x"2000";
    tmp(56254) := x"2000";
    tmp(56255) := x"2800";
    tmp(56256) := x"2000";
    tmp(56257) := x"1800";
    tmp(56258) := x"1800";
    tmp(56259) := x"1800";
    tmp(56260) := x"1800";
    tmp(56261) := x"2000";
    tmp(56262) := x"2800";
    tmp(56263) := x"2800";
    tmp(56264) := x"2800";
    tmp(56265) := x"2800";
    tmp(56266) := x"3000";
    tmp(56267) := x"3800";
    tmp(56268) := x"4000";
    tmp(56269) := x"4000";
    tmp(56270) := x"3800";
    tmp(56271) := x"3800";
    tmp(56272) := x"3800";
    tmp(56273) := x"3800";
    tmp(56274) := x"3000";
    tmp(56275) := x"3000";
    tmp(56276) := x"3000";
    tmp(56277) := x"3000";
    tmp(56278) := x"3000";
    tmp(56279) := x"3820";
    tmp(56280) := x"3020";
    tmp(56281) := x"2000";
    tmp(56282) := x"2000";
    tmp(56283) := x"2820";
    tmp(56284) := x"50a3";
    tmp(56285) := x"6945";
    tmp(56286) := x"7966";
    tmp(56287) := x"8986";
    tmp(56288) := x"8986";
    tmp(56289) := x"8146";
    tmp(56290) := x"8966";
    tmp(56291) := x"aa09";
    tmp(56292) := x"a209";
    tmp(56293) := x"a1e9";
    tmp(56294) := x"7946";
    tmp(56295) := x"c208";
    tmp(56296) := x"3820";
    tmp(56297) := x"5061";
    tmp(56298) := x"dacc";
    tmp(56299) := x"7082";
    tmp(56300) := x"5041";
    tmp(56301) := x"ca29";
    tmp(56302) := x"68a2";
    tmp(56303) := x"88e4";
    tmp(56304) := x"5841";
    tmp(56305) := x"5020";
    tmp(56306) := x"88a2";
    tmp(56307) := x"e28b";
    tmp(56308) := x"4020";
    tmp(56309) := x"8882";
    tmp(56310) := x"d186";
    tmp(56311) := x"e24a";
    tmp(56312) := x"6861";
    tmp(56313) := x"8882";
    tmp(56314) := x"ea6a";
    tmp(56315) := x"90c3";
    tmp(56316) := x"6841";
    tmp(56317) := x"d208";
    tmp(56318) := x"b145";
    tmp(56319) := x"6841";
    tmp(56320) := x"5020";
    tmp(56321) := x"6041";
    tmp(56322) := x"2800";
    tmp(56323) := x"2800";
    tmp(56324) := x"2000";
    tmp(56325) := x"2000";
    tmp(56326) := x"3800";
    tmp(56327) := x"4800";
    tmp(56328) := x"5800";
    tmp(56329) := x"6000";
    tmp(56330) := x"6800";
    tmp(56331) := x"7000";
    tmp(56332) := x"8800";
    tmp(56333) := x"7800";
    tmp(56334) := x"8000";
    tmp(56335) := x"8800";
    tmp(56336) := x"8800";
    tmp(56337) := x"8800";
    tmp(56338) := x"9800";
    tmp(56339) := x"9000";
    tmp(56340) := x"a000";
    tmp(56341) := x"c020";
    tmp(56342) := x"c820";
    tmp(56343) := x"b000";
    tmp(56344) := x"b000";
    tmp(56345) := x"d020";
    tmp(56346) := x"8820";
    tmp(56347) := x"2040";
    tmp(56348) := x"0840";
    tmp(56349) := x"0841";
    tmp(56350) := x"0840";
    tmp(56351) := x"0840";
    tmp(56352) := x"0840";
    tmp(56353) := x"0840";
    tmp(56354) := x"0840";
    tmp(56355) := x"0840";
    tmp(56356) := x"0840";
    tmp(56357) := x"0840";
    tmp(56358) := x"0840";
    tmp(56359) := x"0840";
    tmp(56360) := x"0840";
    tmp(56361) := x"0840";
    tmp(56362) := x"0840";
    tmp(56363) := x"0840";
    tmp(56364) := x"0840";
    tmp(56365) := x"0820";
    tmp(56366) := x"0820";
    tmp(56367) := x"0820";
    tmp(56368) := x"0820";
    tmp(56369) := x"0820";
    tmp(56370) := x"0820";
    tmp(56371) := x"0820";
    tmp(56372) := x"0820";
    tmp(56373) := x"0820";
    tmp(56374) := x"0820";
    tmp(56375) := x"0820";
    tmp(56376) := x"0820";
    tmp(56377) := x"0820";
    tmp(56378) := x"0020";
    tmp(56379) := x"0020";
    tmp(56380) := x"0820";
    tmp(56381) := x"0820";
    tmp(56382) := x"0820";
    tmp(56383) := x"0820";
    tmp(56384) := x"0820";
    tmp(56385) := x"0820";
    tmp(56386) := x"0820";
    tmp(56387) := x"0820";
    tmp(56388) := x"0820";
    tmp(56389) := x"0820";
    tmp(56390) := x"0820";
    tmp(56391) := x"0820";
    tmp(56392) := x"0820";
    tmp(56393) := x"0820";
    tmp(56394) := x"0820";
    tmp(56395) := x"0820";
    tmp(56396) := x"0820";
    tmp(56397) := x"0820";
    tmp(56398) := x"0820";
    tmp(56399) := x"0820";
    tmp(56400) := x"0000";
    tmp(56401) := x"0800";
    tmp(56402) := x"1000";
    tmp(56403) := x"1000";
    tmp(56404) := x"1000";
    tmp(56405) := x"1800";
    tmp(56406) := x"1000";
    tmp(56407) := x"1800";
    tmp(56408) := x"1000";
    tmp(56409) := x"1000";
    tmp(56410) := x"1000";
    tmp(56411) := x"1000";
    tmp(56412) := x"1000";
    tmp(56413) := x"1000";
    tmp(56414) := x"1000";
    tmp(56415) := x"1000";
    tmp(56416) := x"1800";
    tmp(56417) := x"1800";
    tmp(56418) := x"1800";
    tmp(56419) := x"1800";
    tmp(56420) := x"1800";
    tmp(56421) := x"1800";
    tmp(56422) := x"2000";
    tmp(56423) := x"2000";
    tmp(56424) := x"1800";
    tmp(56425) := x"2000";
    tmp(56426) := x"2000";
    tmp(56427) := x"1800";
    tmp(56428) := x"1800";
    tmp(56429) := x"1800";
    tmp(56430) := x"2000";
    tmp(56431) := x"2000";
    tmp(56432) := x"2000";
    tmp(56433) := x"2000";
    tmp(56434) := x"2000";
    tmp(56435) := x"2000";
    tmp(56436) := x"2000";
    tmp(56437) := x"2800";
    tmp(56438) := x"2800";
    tmp(56439) := x"2800";
    tmp(56440) := x"2800";
    tmp(56441) := x"2000";
    tmp(56442) := x"2000";
    tmp(56443) := x"2800";
    tmp(56444) := x"3000";
    tmp(56445) := x"3000";
    tmp(56446) := x"2800";
    tmp(56447) := x"2800";
    tmp(56448) := x"3000";
    tmp(56449) := x"3000";
    tmp(56450) := x"3000";
    tmp(56451) := x"3000";
    tmp(56452) := x"2800";
    tmp(56453) := x"2800";
    tmp(56454) := x"3000";
    tmp(56455) := x"3000";
    tmp(56456) := x"3000";
    tmp(56457) := x"3000";
    tmp(56458) := x"3000";
    tmp(56459) := x"3000";
    tmp(56460) := x"3000";
    tmp(56461) := x"3000";
    tmp(56462) := x"3000";
    tmp(56463) := x"3000";
    tmp(56464) := x"2800";
    tmp(56465) := x"2800";
    tmp(56466) := x"2000";
    tmp(56467) := x"2800";
    tmp(56468) := x"2000";
    tmp(56469) := x"2000";
    tmp(56470) := x"2000";
    tmp(56471) := x"2000";
    tmp(56472) := x"1800";
    tmp(56473) := x"1800";
    tmp(56474) := x"1800";
    tmp(56475) := x"1800";
    tmp(56476) := x"1800";
    tmp(56477) := x"2000";
    tmp(56478) := x"2000";
    tmp(56479) := x"2000";
    tmp(56480) := x"2000";
    tmp(56481) := x"2000";
    tmp(56482) := x"2000";
    tmp(56483) := x"2000";
    tmp(56484) := x"2000";
    tmp(56485) := x"2000";
    tmp(56486) := x"1800";
    tmp(56487) := x"1800";
    tmp(56488) := x"1000";
    tmp(56489) := x"1000";
    tmp(56490) := x"1000";
    tmp(56491) := x"1800";
    tmp(56492) := x"2000";
    tmp(56493) := x"2000";
    tmp(56494) := x"2800";
    tmp(56495) := x"2800";
    tmp(56496) := x"2000";
    tmp(56497) := x"1800";
    tmp(56498) := x"1800";
    tmp(56499) := x"1800";
    tmp(56500) := x"2800";
    tmp(56501) := x"3000";
    tmp(56502) := x"3800";
    tmp(56503) := x"3800";
    tmp(56504) := x"3000";
    tmp(56505) := x"3000";
    tmp(56506) := x"3800";
    tmp(56507) := x"4000";
    tmp(56508) := x"4800";
    tmp(56509) := x"4800";
    tmp(56510) := x"4000";
    tmp(56511) := x"4000";
    tmp(56512) := x"4800";
    tmp(56513) := x"5000";
    tmp(56514) := x"4800";
    tmp(56515) := x"4020";
    tmp(56516) := x"3000";
    tmp(56517) := x"3800";
    tmp(56518) := x"4020";
    tmp(56519) := x"4820";
    tmp(56520) := x"4820";
    tmp(56521) := x"5020";
    tmp(56522) := x"5020";
    tmp(56523) := x"4821";
    tmp(56524) := x"3841";
    tmp(56525) := x"3862";
    tmp(56526) := x"40a2";
    tmp(56527) := x"58e4";
    tmp(56528) := x"58e4";
    tmp(56529) := x"7966";
    tmp(56530) := x"a208";
    tmp(56531) := x"b24a";
    tmp(56532) := x"8987";
    tmp(56533) := x"91a7";
    tmp(56534) := x"9187";
    tmp(56535) := x"70a2";
    tmp(56536) := x"3800";
    tmp(56537) := x"6861";
    tmp(56538) := x"9145";
    tmp(56539) := x"6041";
    tmp(56540) := x"6041";
    tmp(56541) := x"c229";
    tmp(56542) := x"5041";
    tmp(56543) := x"5841";
    tmp(56544) := x"5020";
    tmp(56545) := x"5820";
    tmp(56546) := x"5020";
    tmp(56547) := x"e2ab";
    tmp(56548) := x"a904";
    tmp(56549) := x"6861";
    tmp(56550) := x"b924";
    tmp(56551) := x"90e3";
    tmp(56552) := x"c165";
    tmp(56553) := x"5820";
    tmp(56554) := x"c904";
    tmp(56555) := x"b904";
    tmp(56556) := x"5020";
    tmp(56557) := x"9882";
    tmp(56558) := x"c104";
    tmp(56559) := x"7841";
    tmp(56560) := x"5820";
    tmp(56561) := x"4000";
    tmp(56562) := x"2800";
    tmp(56563) := x"2800";
    tmp(56564) := x"2800";
    tmp(56565) := x"2800";
    tmp(56566) := x"3000";
    tmp(56567) := x"4800";
    tmp(56568) := x"5000";
    tmp(56569) := x"6000";
    tmp(56570) := x"6800";
    tmp(56571) := x"7000";
    tmp(56572) := x"9020";
    tmp(56573) := x"9020";
    tmp(56574) := x"8800";
    tmp(56575) := x"8800";
    tmp(56576) := x"9000";
    tmp(56577) := x"9000";
    tmp(56578) := x"9800";
    tmp(56579) := x"9000";
    tmp(56580) := x"a820";
    tmp(56581) := x"b820";
    tmp(56582) := x"a000";
    tmp(56583) := x"b020";
    tmp(56584) := x"b820";
    tmp(56585) := x"c820";
    tmp(56586) := x"7840";
    tmp(56587) := x"1840";
    tmp(56588) := x"0840";
    tmp(56589) := x"0841";
    tmp(56590) := x"0841";
    tmp(56591) := x"0840";
    tmp(56592) := x"0840";
    tmp(56593) := x"0841";
    tmp(56594) := x"0840";
    tmp(56595) := x"0840";
    tmp(56596) := x"0840";
    tmp(56597) := x"0840";
    tmp(56598) := x"0840";
    tmp(56599) := x"0840";
    tmp(56600) := x"0840";
    tmp(56601) := x"0840";
    tmp(56602) := x"0820";
    tmp(56603) := x"0820";
    tmp(56604) := x"0820";
    tmp(56605) := x"0820";
    tmp(56606) := x"0820";
    tmp(56607) := x"0820";
    tmp(56608) := x"0820";
    tmp(56609) := x"0820";
    tmp(56610) := x"0820";
    tmp(56611) := x"0820";
    tmp(56612) := x"0820";
    tmp(56613) := x"0820";
    tmp(56614) := x"0820";
    tmp(56615) := x"0820";
    tmp(56616) := x"0820";
    tmp(56617) := x"0820";
    tmp(56618) := x"0820";
    tmp(56619) := x"0820";
    tmp(56620) := x"0820";
    tmp(56621) := x"0820";
    tmp(56622) := x"0820";
    tmp(56623) := x"0820";
    tmp(56624) := x"0820";
    tmp(56625) := x"0820";
    tmp(56626) := x"0820";
    tmp(56627) := x"0820";
    tmp(56628) := x"0820";
    tmp(56629) := x"0820";
    tmp(56630) := x"0820";
    tmp(56631) := x"0820";
    tmp(56632) := x"0820";
    tmp(56633) := x"0820";
    tmp(56634) := x"0820";
    tmp(56635) := x"0840";
    tmp(56636) := x"0820";
    tmp(56637) := x"0820";
    tmp(56638) := x"0820";
    tmp(56639) := x"0820";
    tmp(56640) := x"0000";
    tmp(56641) := x"1000";
    tmp(56642) := x"1000";
    tmp(56643) := x"1000";
    tmp(56644) := x"1000";
    tmp(56645) := x"1000";
    tmp(56646) := x"1000";
    tmp(56647) := x"1000";
    tmp(56648) := x"1000";
    tmp(56649) := x"0800";
    tmp(56650) := x"0800";
    tmp(56651) := x"1000";
    tmp(56652) := x"1000";
    tmp(56653) := x"1800";
    tmp(56654) := x"1800";
    tmp(56655) := x"1800";
    tmp(56656) := x"1800";
    tmp(56657) := x"1800";
    tmp(56658) := x"1800";
    tmp(56659) := x"1800";
    tmp(56660) := x"1800";
    tmp(56661) := x"1800";
    tmp(56662) := x"1000";
    tmp(56663) := x"1000";
    tmp(56664) := x"1000";
    tmp(56665) := x"1800";
    tmp(56666) := x"1800";
    tmp(56667) := x"1800";
    tmp(56668) := x"1800";
    tmp(56669) := x"2000";
    tmp(56670) := x"2000";
    tmp(56671) := x"2000";
    tmp(56672) := x"2000";
    tmp(56673) := x"2000";
    tmp(56674) := x"2000";
    tmp(56675) := x"2000";
    tmp(56676) := x"2000";
    tmp(56677) := x"2000";
    tmp(56678) := x"2000";
    tmp(56679) := x"2000";
    tmp(56680) := x"2800";
    tmp(56681) := x"2800";
    tmp(56682) := x"2800";
    tmp(56683) := x"2800";
    tmp(56684) := x"3000";
    tmp(56685) := x"3000";
    tmp(56686) := x"2800";
    tmp(56687) := x"2800";
    tmp(56688) := x"2000";
    tmp(56689) := x"2000";
    tmp(56690) := x"2800";
    tmp(56691) := x"2800";
    tmp(56692) := x"2800";
    tmp(56693) := x"2800";
    tmp(56694) := x"2800";
    tmp(56695) := x"3000";
    tmp(56696) := x"3000";
    tmp(56697) := x"3000";
    tmp(56698) := x"3000";
    tmp(56699) := x"3000";
    tmp(56700) := x"3000";
    tmp(56701) := x"3000";
    tmp(56702) := x"3000";
    tmp(56703) := x"3000";
    tmp(56704) := x"2800";
    tmp(56705) := x"2000";
    tmp(56706) := x"2000";
    tmp(56707) := x"2000";
    tmp(56708) := x"2000";
    tmp(56709) := x"2000";
    tmp(56710) := x"2000";
    tmp(56711) := x"2000";
    tmp(56712) := x"2000";
    tmp(56713) := x"2000";
    tmp(56714) := x"2000";
    tmp(56715) := x"1800";
    tmp(56716) := x"1800";
    tmp(56717) := x"1800";
    tmp(56718) := x"2000";
    tmp(56719) := x"2000";
    tmp(56720) := x"2000";
    tmp(56721) := x"2000";
    tmp(56722) := x"2000";
    tmp(56723) := x"2000";
    tmp(56724) := x"2000";
    tmp(56725) := x"2000";
    tmp(56726) := x"2000";
    tmp(56727) := x"1800";
    tmp(56728) := x"1000";
    tmp(56729) := x"1000";
    tmp(56730) := x"1000";
    tmp(56731) := x"1000";
    tmp(56732) := x"1800";
    tmp(56733) := x"2000";
    tmp(56734) := x"2800";
    tmp(56735) := x"2800";
    tmp(56736) := x"2000";
    tmp(56737) := x"2000";
    tmp(56738) := x"2800";
    tmp(56739) := x"3000";
    tmp(56740) := x"3000";
    tmp(56741) := x"3800";
    tmp(56742) := x"3800";
    tmp(56743) := x"3800";
    tmp(56744) := x"3000";
    tmp(56745) := x"3000";
    tmp(56746) := x"3800";
    tmp(56747) := x"4000";
    tmp(56748) := x"4000";
    tmp(56749) := x"4800";
    tmp(56750) := x"4000";
    tmp(56751) := x"4000";
    tmp(56752) := x"4800";
    tmp(56753) := x"5000";
    tmp(56754) := x"4800";
    tmp(56755) := x"4000";
    tmp(56756) := x"4000";
    tmp(56757) := x"4800";
    tmp(56758) := x"5000";
    tmp(56759) := x"5020";
    tmp(56760) := x"5820";
    tmp(56761) := x"6820";
    tmp(56762) := x"6820";
    tmp(56763) := x"7021";
    tmp(56764) := x"6041";
    tmp(56765) := x"5061";
    tmp(56766) := x"48a2";
    tmp(56767) := x"60e3";
    tmp(56768) := x"68e3";
    tmp(56769) := x"58a2";
    tmp(56770) := x"8125";
    tmp(56771) := x"8966";
    tmp(56772) := x"8986";
    tmp(56773) := x"9187";
    tmp(56774) := x"b9e8";
    tmp(56775) := x"5021";
    tmp(56776) := x"5020";
    tmp(56777) := x"6041";
    tmp(56778) := x"78a2";
    tmp(56779) := x"4820";
    tmp(56780) := x"5841";
    tmp(56781) := x"80e3";
    tmp(56782) := x"4820";
    tmp(56783) := x"4800";
    tmp(56784) := x"5020";
    tmp(56785) := x"6820";
    tmp(56786) := x"4800";
    tmp(56787) := x"8861";
    tmp(56788) := x"d9c6";
    tmp(56789) := x"88a2";
    tmp(56790) := x"9082";
    tmp(56791) := x"6020";
    tmp(56792) := x"9061";
    tmp(56793) := x"5800";
    tmp(56794) := x"7021";
    tmp(56795) := x"c124";
    tmp(56796) := x"7841";
    tmp(56797) := x"6020";
    tmp(56798) := x"7820";
    tmp(56799) := x"6820";
    tmp(56800) := x"6020";
    tmp(56801) := x"4000";
    tmp(56802) := x"3000";
    tmp(56803) := x"3000";
    tmp(56804) := x"3000";
    tmp(56805) := x"3000";
    tmp(56806) := x"3800";
    tmp(56807) := x"4800";
    tmp(56808) := x"5000";
    tmp(56809) := x"6000";
    tmp(56810) := x"6800";
    tmp(56811) := x"7000";
    tmp(56812) := x"8000";
    tmp(56813) := x"8000";
    tmp(56814) := x"8000";
    tmp(56815) := x"9000";
    tmp(56816) := x"9000";
    tmp(56817) := x"a000";
    tmp(56818) := x"a000";
    tmp(56819) := x"9800";
    tmp(56820) := x"a800";
    tmp(56821) := x"9000";
    tmp(56822) := x"a800";
    tmp(56823) := x"c820";
    tmp(56824) := x"d820";
    tmp(56825) := x"c820";
    tmp(56826) := x"7860";
    tmp(56827) := x"1840";
    tmp(56828) := x"0841";
    tmp(56829) := x"0841";
    tmp(56830) := x"0841";
    tmp(56831) := x"0840";
    tmp(56832) := x"0840";
    tmp(56833) := x"0840";
    tmp(56834) := x"0840";
    tmp(56835) := x"0840";
    tmp(56836) := x"0840";
    tmp(56837) := x"0840";
    tmp(56838) := x"0840";
    tmp(56839) := x"0840";
    tmp(56840) := x"0840";
    tmp(56841) := x"0840";
    tmp(56842) := x"0820";
    tmp(56843) := x"0820";
    tmp(56844) := x"0820";
    tmp(56845) := x"0840";
    tmp(56846) := x"0840";
    tmp(56847) := x"0840";
    tmp(56848) := x"0840";
    tmp(56849) := x"0840";
    tmp(56850) := x"0840";
    tmp(56851) := x"0840";
    tmp(56852) := x"0840";
    tmp(56853) := x"0840";
    tmp(56854) := x"0840";
    tmp(56855) := x"0840";
    tmp(56856) := x"0841";
    tmp(56857) := x"0841";
    tmp(56858) := x"0841";
    tmp(56859) := x"0841";
    tmp(56860) := x"0840";
    tmp(56861) := x"0840";
    tmp(56862) := x"0840";
    tmp(56863) := x"0840";
    tmp(56864) := x"0840";
    tmp(56865) := x"0840";
    tmp(56866) := x"0840";
    tmp(56867) := x"0840";
    tmp(56868) := x"0840";
    tmp(56869) := x"0840";
    tmp(56870) := x"0840";
    tmp(56871) := x"0840";
    tmp(56872) := x"0840";
    tmp(56873) := x"0840";
    tmp(56874) := x"0840";
    tmp(56875) := x"0840";
    tmp(56876) := x"0840";
    tmp(56877) := x"0840";
    tmp(56878) := x"0840";
    tmp(56879) := x"0820";
    tmp(56880) := x"0000";
    tmp(56881) := x"0800";
    tmp(56882) := x"1000";
    tmp(56883) := x"1000";
    tmp(56884) := x"1000";
    tmp(56885) := x"1000";
    tmp(56886) := x"1000";
    tmp(56887) := x"0800";
    tmp(56888) := x"0800";
    tmp(56889) := x"1000";
    tmp(56890) := x"1000";
    tmp(56891) := x"1000";
    tmp(56892) := x"1000";
    tmp(56893) := x"1800";
    tmp(56894) := x"1800";
    tmp(56895) := x"1800";
    tmp(56896) := x"1800";
    tmp(56897) := x"1800";
    tmp(56898) := x"1800";
    tmp(56899) := x"1000";
    tmp(56900) := x"1000";
    tmp(56901) := x"1000";
    tmp(56902) := x"1000";
    tmp(56903) := x"1000";
    tmp(56904) := x"1000";
    tmp(56905) := x"1800";
    tmp(56906) := x"1800";
    tmp(56907) := x"1800";
    tmp(56908) := x"2000";
    tmp(56909) := x"2000";
    tmp(56910) := x"2000";
    tmp(56911) := x"2000";
    tmp(56912) := x"2000";
    tmp(56913) := x"1800";
    tmp(56914) := x"1800";
    tmp(56915) := x"1800";
    tmp(56916) := x"2000";
    tmp(56917) := x"2000";
    tmp(56918) := x"2000";
    tmp(56919) := x"2000";
    tmp(56920) := x"2800";
    tmp(56921) := x"2800";
    tmp(56922) := x"2800";
    tmp(56923) := x"2800";
    tmp(56924) := x"2800";
    tmp(56925) := x"2800";
    tmp(56926) := x"2800";
    tmp(56927) := x"2800";
    tmp(56928) := x"2800";
    tmp(56929) := x"2800";
    tmp(56930) := x"2800";
    tmp(56931) := x"2800";
    tmp(56932) := x"2800";
    tmp(56933) := x"2800";
    tmp(56934) := x"3000";
    tmp(56935) := x"3000";
    tmp(56936) := x"3000";
    tmp(56937) := x"3000";
    tmp(56938) := x"3000";
    tmp(56939) := x"3000";
    tmp(56940) := x"3000";
    tmp(56941) := x"3000";
    tmp(56942) := x"3000";
    tmp(56943) := x"3000";
    tmp(56944) := x"2800";
    tmp(56945) := x"2800";
    tmp(56946) := x"2000";
    tmp(56947) := x"1800";
    tmp(56948) := x"2000";
    tmp(56949) := x"2000";
    tmp(56950) := x"2800";
    tmp(56951) := x"2800";
    tmp(56952) := x"2800";
    tmp(56953) := x"2800";
    tmp(56954) := x"2000";
    tmp(56955) := x"2000";
    tmp(56956) := x"2000";
    tmp(56957) := x"2000";
    tmp(56958) := x"1800";
    tmp(56959) := x"2000";
    tmp(56960) := x"2000";
    tmp(56961) := x"2800";
    tmp(56962) := x"2800";
    tmp(56963) := x"2800";
    tmp(56964) := x"2000";
    tmp(56965) := x"2000";
    tmp(56966) := x"1800";
    tmp(56967) := x"1800";
    tmp(56968) := x"1000";
    tmp(56969) := x"1000";
    tmp(56970) := x"1000";
    tmp(56971) := x"1000";
    tmp(56972) := x"1800";
    tmp(56973) := x"1800";
    tmp(56974) := x"2000";
    tmp(56975) := x"2000";
    tmp(56976) := x"2000";
    tmp(56977) := x"2000";
    tmp(56978) := x"2800";
    tmp(56979) := x"2800";
    tmp(56980) := x"3000";
    tmp(56981) := x"3800";
    tmp(56982) := x"3800";
    tmp(56983) := x"3800";
    tmp(56984) := x"3800";
    tmp(56985) := x"3000";
    tmp(56986) := x"3800";
    tmp(56987) := x"4000";
    tmp(56988) := x"4000";
    tmp(56989) := x"4000";
    tmp(56990) := x"4800";
    tmp(56991) := x"4000";
    tmp(56992) := x"4000";
    tmp(56993) := x"5000";
    tmp(56994) := x"4800";
    tmp(56995) := x"4000";
    tmp(56996) := x"4000";
    tmp(56997) := x"4000";
    tmp(56998) := x"5000";
    tmp(56999) := x"5000";
    tmp(57000) := x"5000";
    tmp(57001) := x"6000";
    tmp(57002) := x"6820";
    tmp(57003) := x"6820";
    tmp(57004) := x"6020";
    tmp(57005) := x"4820";
    tmp(57006) := x"4021";
    tmp(57007) := x"3820";
    tmp(57008) := x"3820";
    tmp(57009) := x"4020";
    tmp(57010) := x"4820";
    tmp(57011) := x"6882";
    tmp(57012) := x"7904";
    tmp(57013) := x"70e3";
    tmp(57014) := x"6882";
    tmp(57015) := x"5020";
    tmp(57016) := x"5820";
    tmp(57017) := x"7061";
    tmp(57018) := x"80a2";
    tmp(57019) := x"3800";
    tmp(57020) := x"6841";
    tmp(57021) := x"90e4";
    tmp(57022) := x"4020";
    tmp(57023) := x"4800";
    tmp(57024) := x"5820";
    tmp(57025) := x"8881";
    tmp(57026) := x"6020";
    tmp(57027) := x"5000";
    tmp(57028) := x"a8a2";
    tmp(57029) := x"7841";
    tmp(57030) := x"7841";
    tmp(57031) := x"7020";
    tmp(57032) := x"7020";
    tmp(57033) := x"7020";
    tmp(57034) := x"6000";
    tmp(57035) := x"8861";
    tmp(57036) := x"9881";
    tmp(57037) := x"7820";
    tmp(57038) := x"6820";
    tmp(57039) := x"6820";
    tmp(57040) := x"6020";
    tmp(57041) := x"4000";
    tmp(57042) := x"3000";
    tmp(57043) := x"3800";
    tmp(57044) := x"3000";
    tmp(57045) := x"3000";
    tmp(57046) := x"3800";
    tmp(57047) := x"4800";
    tmp(57048) := x"5800";
    tmp(57049) := x"6000";
    tmp(57050) := x"6000";
    tmp(57051) := x"7800";
    tmp(57052) := x"8000";
    tmp(57053) := x"8000";
    tmp(57054) := x"8800";
    tmp(57055) := x"9800";
    tmp(57056) := x"9800";
    tmp(57057) := x"a000";
    tmp(57058) := x"a000";
    tmp(57059) := x"a000";
    tmp(57060) := x"a800";
    tmp(57061) := x"9800";
    tmp(57062) := x"b820";
    tmp(57063) := x"d020";
    tmp(57064) := x"f840";
    tmp(57065) := x"e860";
    tmp(57066) := x"6881";
    tmp(57067) := x"1040";
    tmp(57068) := x"0841";
    tmp(57069) := x"0841";
    tmp(57070) := x"0840";
    tmp(57071) := x"0841";
    tmp(57072) := x"0840";
    tmp(57073) := x"0840";
    tmp(57074) := x"0840";
    tmp(57075) := x"0840";
    tmp(57076) := x"0840";
    tmp(57077) := x"0840";
    tmp(57078) := x"0840";
    tmp(57079) := x"0840";
    tmp(57080) := x"0840";
    tmp(57081) := x"0840";
    tmp(57082) := x"0840";
    tmp(57083) := x"0840";
    tmp(57084) := x"0840";
    tmp(57085) := x"0841";
    tmp(57086) := x"0841";
    tmp(57087) := x"0841";
    tmp(57088) := x"0841";
    tmp(57089) := x"0861";
    tmp(57090) := x"0841";
    tmp(57091) := x"0841";
    tmp(57092) := x"0841";
    tmp(57093) := x"0861";
    tmp(57094) := x"0861";
    tmp(57095) := x"0861";
    tmp(57096) := x"0861";
    tmp(57097) := x"0861";
    tmp(57098) := x"0861";
    tmp(57099) := x"0861";
    tmp(57100) := x"0861";
    tmp(57101) := x"0861";
    tmp(57102) := x"0861";
    tmp(57103) := x"0861";
    tmp(57104) := x"0841";
    tmp(57105) := x"0841";
    tmp(57106) := x"0841";
    tmp(57107) := x"0841";
    tmp(57108) := x"0840";
    tmp(57109) := x"0840";
    tmp(57110) := x"0840";
    tmp(57111) := x"0840";
    tmp(57112) := x"0841";
    tmp(57113) := x"0841";
    tmp(57114) := x"0840";
    tmp(57115) := x"0841";
    tmp(57116) := x"0840";
    tmp(57117) := x"0840";
    tmp(57118) := x"0840";
    tmp(57119) := x"0840";
    tmp(57120) := x"0000";
    tmp(57121) := x"1000";
    tmp(57122) := x"1000";
    tmp(57123) := x"1000";
    tmp(57124) := x"0800";
    tmp(57125) := x"0800";
    tmp(57126) := x"0800";
    tmp(57127) := x"0800";
    tmp(57128) := x"1000";
    tmp(57129) := x"1000";
    tmp(57130) := x"1000";
    tmp(57131) := x"1000";
    tmp(57132) := x"1000";
    tmp(57133) := x"1800";
    tmp(57134) := x"1800";
    tmp(57135) := x"1800";
    tmp(57136) := x"1800";
    tmp(57137) := x"1800";
    tmp(57138) := x"1000";
    tmp(57139) := x"1000";
    tmp(57140) := x"1000";
    tmp(57141) := x"1000";
    tmp(57142) := x"1000";
    tmp(57143) := x"1000";
    tmp(57144) := x"1000";
    tmp(57145) := x"1800";
    tmp(57146) := x"1800";
    tmp(57147) := x"1800";
    tmp(57148) := x"2000";
    tmp(57149) := x"2000";
    tmp(57150) := x"2000";
    tmp(57151) := x"2000";
    tmp(57152) := x"1800";
    tmp(57153) := x"1800";
    tmp(57154) := x"1800";
    tmp(57155) := x"1800";
    tmp(57156) := x"1800";
    tmp(57157) := x"2000";
    tmp(57158) := x"2000";
    tmp(57159) := x"2000";
    tmp(57160) := x"2000";
    tmp(57161) := x"2800";
    tmp(57162) := x"2800";
    tmp(57163) := x"2800";
    tmp(57164) := x"2800";
    tmp(57165) := x"2800";
    tmp(57166) := x"2800";
    tmp(57167) := x"3000";
    tmp(57168) := x"2800";
    tmp(57169) := x"2800";
    tmp(57170) := x"2800";
    tmp(57171) := x"2800";
    tmp(57172) := x"2800";
    tmp(57173) := x"2800";
    tmp(57174) := x"2800";
    tmp(57175) := x"2800";
    tmp(57176) := x"2800";
    tmp(57177) := x"2800";
    tmp(57178) := x"2800";
    tmp(57179) := x"2800";
    tmp(57180) := x"2800";
    tmp(57181) := x"2800";
    tmp(57182) := x"2800";
    tmp(57183) := x"2800";
    tmp(57184) := x"2800";
    tmp(57185) := x"2000";
    tmp(57186) := x"2000";
    tmp(57187) := x"1800";
    tmp(57188) := x"2000";
    tmp(57189) := x"2800";
    tmp(57190) := x"2800";
    tmp(57191) := x"2800";
    tmp(57192) := x"2800";
    tmp(57193) := x"2800";
    tmp(57194) := x"2800";
    tmp(57195) := x"2000";
    tmp(57196) := x"2000";
    tmp(57197) := x"2000";
    tmp(57198) := x"2000";
    tmp(57199) := x"2000";
    tmp(57200) := x"2000";
    tmp(57201) := x"2000";
    tmp(57202) := x"2000";
    tmp(57203) := x"2000";
    tmp(57204) := x"2000";
    tmp(57205) := x"2000";
    tmp(57206) := x"2000";
    tmp(57207) := x"1800";
    tmp(57208) := x"1800";
    tmp(57209) := x"1000";
    tmp(57210) := x"1000";
    tmp(57211) := x"1000";
    tmp(57212) := x"1000";
    tmp(57213) := x"1800";
    tmp(57214) := x"2000";
    tmp(57215) := x"1800";
    tmp(57216) := x"1800";
    tmp(57217) := x"1000";
    tmp(57218) := x"1000";
    tmp(57219) := x"1000";
    tmp(57220) := x"2000";
    tmp(57221) := x"3000";
    tmp(57222) := x"3800";
    tmp(57223) := x"3800";
    tmp(57224) := x"3800";
    tmp(57225) := x"3800";
    tmp(57226) := x"3800";
    tmp(57227) := x"3800";
    tmp(57228) := x"3800";
    tmp(57229) := x"4000";
    tmp(57230) := x"4800";
    tmp(57231) := x"4000";
    tmp(57232) := x"4000";
    tmp(57233) := x"4000";
    tmp(57234) := x"5000";
    tmp(57235) := x"5000";
    tmp(57236) := x"4000";
    tmp(57237) := x"4800";
    tmp(57238) := x"4800";
    tmp(57239) := x"5000";
    tmp(57240) := x"5800";
    tmp(57241) := x"5800";
    tmp(57242) := x"5800";
    tmp(57243) := x"5800";
    tmp(57244) := x"5000";
    tmp(57245) := x"3800";
    tmp(57246) := x"4000";
    tmp(57247) := x"4800";
    tmp(57248) := x"5820";
    tmp(57249) := x"6820";
    tmp(57250) := x"7820";
    tmp(57251) := x"7841";
    tmp(57252) := x"6861";
    tmp(57253) := x"5841";
    tmp(57254) := x"4820";
    tmp(57255) := x"5820";
    tmp(57256) := x"6020";
    tmp(57257) := x"7061";
    tmp(57258) := x"7881";
    tmp(57259) := x"4800";
    tmp(57260) := x"7041";
    tmp(57261) := x"80a2";
    tmp(57262) := x"4820";
    tmp(57263) := x"4800";
    tmp(57264) := x"5820";
    tmp(57265) := x"7041";
    tmp(57266) := x"5820";
    tmp(57267) := x"5800";
    tmp(57268) := x"6020";
    tmp(57269) := x"8020";
    tmp(57270) := x"7020";
    tmp(57271) := x"6820";
    tmp(57272) := x"7000";
    tmp(57273) := x"7820";
    tmp(57274) := x"6800";
    tmp(57275) := x"6000";
    tmp(57276) := x"7820";
    tmp(57277) := x"8020";
    tmp(57278) := x"7820";
    tmp(57279) := x"8041";
    tmp(57280) := x"6820";
    tmp(57281) := x"5000";
    tmp(57282) := x"3800";
    tmp(57283) := x"3800";
    tmp(57284) := x"3800";
    tmp(57285) := x"3800";
    tmp(57286) := x"4000";
    tmp(57287) := x"5000";
    tmp(57288) := x"6000";
    tmp(57289) := x"6000";
    tmp(57290) := x"6000";
    tmp(57291) := x"7800";
    tmp(57292) := x"9000";
    tmp(57293) := x"9800";
    tmp(57294) := x"9800";
    tmp(57295) := x"9000";
    tmp(57296) := x"9800";
    tmp(57297) := x"a000";
    tmp(57298) := x"a000";
    tmp(57299) := x"a800";
    tmp(57300) := x"b020";
    tmp(57301) := x"b020";
    tmp(57302) := x"b820";
    tmp(57303) := x"d820";
    tmp(57304) := x"f860";
    tmp(57305) := x"c060";
    tmp(57306) := x"4061";
    tmp(57307) := x"1040";
    tmp(57308) := x"0841";
    tmp(57309) := x"0841";
    tmp(57310) := x"0840";
    tmp(57311) := x"0840";
    tmp(57312) := x"0840";
    tmp(57313) := x"0840";
    tmp(57314) := x"0840";
    tmp(57315) := x"0840";
    tmp(57316) := x"0840";
    tmp(57317) := x"0840";
    tmp(57318) := x"0840";
    tmp(57319) := x"0840";
    tmp(57320) := x"0841";
    tmp(57321) := x"0841";
    tmp(57322) := x"0841";
    tmp(57323) := x"0841";
    tmp(57324) := x"0861";
    tmp(57325) := x"0861";
    tmp(57326) := x"0861";
    tmp(57327) := x"0861";
    tmp(57328) := x"0861";
    tmp(57329) := x"0861";
    tmp(57330) := x"1061";
    tmp(57331) := x"1081";
    tmp(57332) := x"1081";
    tmp(57333) := x"1081";
    tmp(57334) := x"1082";
    tmp(57335) := x"10a2";
    tmp(57336) := x"10a2";
    tmp(57337) := x"1082";
    tmp(57338) := x"10a2";
    tmp(57339) := x"1082";
    tmp(57340) := x"1081";
    tmp(57341) := x"1081";
    tmp(57342) := x"1061";
    tmp(57343) := x"1061";
    tmp(57344) := x"1061";
    tmp(57345) := x"0861";
    tmp(57346) := x"0861";
    tmp(57347) := x"0861";
    tmp(57348) := x"0841";
    tmp(57349) := x"0841";
    tmp(57350) := x"0841";
    tmp(57351) := x"0841";
    tmp(57352) := x"0841";
    tmp(57353) := x"0841";
    tmp(57354) := x"0841";
    tmp(57355) := x"0841";
    tmp(57356) := x"0841";
    tmp(57357) := x"0841";
    tmp(57358) := x"0840";
    tmp(57359) := x"0840";
    tmp(57360) := x"0000";
    tmp(57361) := x"1000";
    tmp(57362) := x"0800";
    tmp(57363) := x"0800";
    tmp(57364) := x"0800";
    tmp(57365) := x"0800";
    tmp(57366) := x"0800";
    tmp(57367) := x"0800";
    tmp(57368) := x"0800";
    tmp(57369) := x"0800";
    tmp(57370) := x"1000";
    tmp(57371) := x"1000";
    tmp(57372) := x"1000";
    tmp(57373) := x"1000";
    tmp(57374) := x"1000";
    tmp(57375) := x"1000";
    tmp(57376) := x"1000";
    tmp(57377) := x"1000";
    tmp(57378) := x"1000";
    tmp(57379) := x"1000";
    tmp(57380) := x"1000";
    tmp(57381) := x"1000";
    tmp(57382) := x"1000";
    tmp(57383) := x"1000";
    tmp(57384) := x"1000";
    tmp(57385) := x"1800";
    tmp(57386) := x"1800";
    tmp(57387) := x"1800";
    tmp(57388) := x"2000";
    tmp(57389) := x"2000";
    tmp(57390) := x"2000";
    tmp(57391) := x"1800";
    tmp(57392) := x"1800";
    tmp(57393) := x"1800";
    tmp(57394) := x"1800";
    tmp(57395) := x"1800";
    tmp(57396) := x"1800";
    tmp(57397) := x"1800";
    tmp(57398) := x"2000";
    tmp(57399) := x"2000";
    tmp(57400) := x"2000";
    tmp(57401) := x"2000";
    tmp(57402) := x"2000";
    tmp(57403) := x"2000";
    tmp(57404) := x"2800";
    tmp(57405) := x"2800";
    tmp(57406) := x"2800";
    tmp(57407) := x"2800";
    tmp(57408) := x"2800";
    tmp(57409) := x"2800";
    tmp(57410) := x"2800";
    tmp(57411) := x"2800";
    tmp(57412) := x"2800";
    tmp(57413) := x"3000";
    tmp(57414) := x"2800";
    tmp(57415) := x"2800";
    tmp(57416) := x"2800";
    tmp(57417) := x"2800";
    tmp(57418) := x"2800";
    tmp(57419) := x"2800";
    tmp(57420) := x"2800";
    tmp(57421) := x"2800";
    tmp(57422) := x"2800";
    tmp(57423) := x"2800";
    tmp(57424) := x"2800";
    tmp(57425) := x"2800";
    tmp(57426) := x"2800";
    tmp(57427) := x"2000";
    tmp(57428) := x"2000";
    tmp(57429) := x"2000";
    tmp(57430) := x"1800";
    tmp(57431) := x"2000";
    tmp(57432) := x"1800";
    tmp(57433) := x"1800";
    tmp(57434) := x"1800";
    tmp(57435) := x"1800";
    tmp(57436) := x"1800";
    tmp(57437) := x"1800";
    tmp(57438) := x"1800";
    tmp(57439) := x"2000";
    tmp(57440) := x"2000";
    tmp(57441) := x"2000";
    tmp(57442) := x"2000";
    tmp(57443) := x"2000";
    tmp(57444) := x"2800";
    tmp(57445) := x"2800";
    tmp(57446) := x"2000";
    tmp(57447) := x"1800";
    tmp(57448) := x"1800";
    tmp(57449) := x"1800";
    tmp(57450) := x"1800";
    tmp(57451) := x"1000";
    tmp(57452) := x"1000";
    tmp(57453) := x"1000";
    tmp(57454) := x"1800";
    tmp(57455) := x"1800";
    tmp(57456) := x"1800";
    tmp(57457) := x"1000";
    tmp(57458) := x"1000";
    tmp(57459) := x"1000";
    tmp(57460) := x"1800";
    tmp(57461) := x"2800";
    tmp(57462) := x"3000";
    tmp(57463) := x"3000";
    tmp(57464) := x"3800";
    tmp(57465) := x"4000";
    tmp(57466) := x"3800";
    tmp(57467) := x"3800";
    tmp(57468) := x"3800";
    tmp(57469) := x"3800";
    tmp(57470) := x"3800";
    tmp(57471) := x"3800";
    tmp(57472) := x"4000";
    tmp(57473) := x"4800";
    tmp(57474) := x"5000";
    tmp(57475) := x"5800";
    tmp(57476) := x"4800";
    tmp(57477) := x"5000";
    tmp(57478) := x"4800";
    tmp(57479) := x"5000";
    tmp(57480) := x"5000";
    tmp(57481) := x"5000";
    tmp(57482) := x"5000";
    tmp(57483) := x"5000";
    tmp(57484) := x"5000";
    tmp(57485) := x"4000";
    tmp(57486) := x"4000";
    tmp(57487) := x"4800";
    tmp(57488) := x"5000";
    tmp(57489) := x"5000";
    tmp(57490) := x"5000";
    tmp(57491) := x"5800";
    tmp(57492) := x"4800";
    tmp(57493) := x"4000";
    tmp(57494) := x"5000";
    tmp(57495) := x"5800";
    tmp(57496) := x"5800";
    tmp(57497) := x"6820";
    tmp(57498) := x"7041";
    tmp(57499) := x"6020";
    tmp(57500) := x"7840";
    tmp(57501) := x"7041";
    tmp(57502) := x"4800";
    tmp(57503) := x"4800";
    tmp(57504) := x"5000";
    tmp(57505) := x"5800";
    tmp(57506) := x"5800";
    tmp(57507) := x"5800";
    tmp(57508) := x"6820";
    tmp(57509) := x"7020";
    tmp(57510) := x"7820";
    tmp(57511) := x"6800";
    tmp(57512) := x"6800";
    tmp(57513) := x"7020";
    tmp(57514) := x"7820";
    tmp(57515) := x"6800";
    tmp(57516) := x"7000";
    tmp(57517) := x"8820";
    tmp(57518) := x"8820";
    tmp(57519) := x"7841";
    tmp(57520) := x"5820";
    tmp(57521) := x"6020";
    tmp(57522) := x"4800";
    tmp(57523) := x"3800";
    tmp(57524) := x"3800";
    tmp(57525) := x"4000";
    tmp(57526) := x"4800";
    tmp(57527) := x"5800";
    tmp(57528) := x"5800";
    tmp(57529) := x"6000";
    tmp(57530) := x"7000";
    tmp(57531) := x"9020";
    tmp(57532) := x"a020";
    tmp(57533) := x"b020";
    tmp(57534) := x"a800";
    tmp(57535) := x"a000";
    tmp(57536) := x"a800";
    tmp(57537) := x"a000";
    tmp(57538) := x"9800";
    tmp(57539) := x"b820";
    tmp(57540) := x"c020";
    tmp(57541) := x"b020";
    tmp(57542) := x"c820";
    tmp(57543) := x"d840";
    tmp(57544) := x"f861";
    tmp(57545) := x"8840";
    tmp(57546) := x"1840";
    tmp(57547) := x"0840";
    tmp(57548) := x"0841";
    tmp(57549) := x"0841";
    tmp(57550) := x"0840";
    tmp(57551) := x"0840";
    tmp(57552) := x"0840";
    tmp(57553) := x"0840";
    tmp(57554) := x"0840";
    tmp(57555) := x"0840";
    tmp(57556) := x"0840";
    tmp(57557) := x"0840";
    tmp(57558) := x"0841";
    tmp(57559) := x"0841";
    tmp(57560) := x"0841";
    tmp(57561) := x"0861";
    tmp(57562) := x"0861";
    tmp(57563) := x"1061";
    tmp(57564) := x"1061";
    tmp(57565) := x"1061";
    tmp(57566) := x"1081";
    tmp(57567) := x"1081";
    tmp(57568) := x"1082";
    tmp(57569) := x"1082";
    tmp(57570) := x"10a2";
    tmp(57571) := x"10a2";
    tmp(57572) := x"10a2";
    tmp(57573) := x"10c2";
    tmp(57574) := x"10a3";
    tmp(57575) := x"10c3";
    tmp(57576) := x"18c3";
    tmp(57577) := x"18c3";
    tmp(57578) := x"18c3";
    tmp(57579) := x"10c3";
    tmp(57580) := x"10a2";
    tmp(57581) := x"10a2";
    tmp(57582) := x"10a2";
    tmp(57583) := x"10a2";
    tmp(57584) := x"1081";
    tmp(57585) := x"1081";
    tmp(57586) := x"1061";
    tmp(57587) := x"1061";
    tmp(57588) := x"0861";
    tmp(57589) := x"0861";
    tmp(57590) := x"0841";
    tmp(57591) := x"0841";
    tmp(57592) := x"0841";
    tmp(57593) := x"0841";
    tmp(57594) := x"0841";
    tmp(57595) := x"0841";
    tmp(57596) := x"0841";
    tmp(57597) := x"0841";
    tmp(57598) := x"0841";
    tmp(57599) := x"0840";
    tmp(57600) := x"0000";
    tmp(57601) := x"0800";
    tmp(57602) := x"0800";
    tmp(57603) := x"0800";
    tmp(57604) := x"0800";
    tmp(57605) := x"0800";
    tmp(57606) := x"0800";
    tmp(57607) := x"0800";
    tmp(57608) := x"0800";
    tmp(57609) := x"0800";
    tmp(57610) := x"0800";
    tmp(57611) := x"1000";
    tmp(57612) := x"1000";
    tmp(57613) := x"1000";
    tmp(57614) := x"1000";
    tmp(57615) := x"1000";
    tmp(57616) := x"1000";
    tmp(57617) := x"1000";
    tmp(57618) := x"1000";
    tmp(57619) := x"1000";
    tmp(57620) := x"1000";
    tmp(57621) := x"1000";
    tmp(57622) := x"1000";
    tmp(57623) := x"1000";
    tmp(57624) := x"1000";
    tmp(57625) := x"1800";
    tmp(57626) := x"1800";
    tmp(57627) := x"1800";
    tmp(57628) := x"1800";
    tmp(57629) := x"1800";
    tmp(57630) := x"1800";
    tmp(57631) := x"1800";
    tmp(57632) := x"1800";
    tmp(57633) := x"1800";
    tmp(57634) := x"2000";
    tmp(57635) := x"2000";
    tmp(57636) := x"2000";
    tmp(57637) := x"2000";
    tmp(57638) := x"2000";
    tmp(57639) := x"2000";
    tmp(57640) := x"2000";
    tmp(57641) := x"2000";
    tmp(57642) := x"2000";
    tmp(57643) := x"2000";
    tmp(57644) := x"2800";
    tmp(57645) := x"2800";
    tmp(57646) := x"2800";
    tmp(57647) := x"2800";
    tmp(57648) := x"2800";
    tmp(57649) := x"2800";
    tmp(57650) := x"2800";
    tmp(57651) := x"2800";
    tmp(57652) := x"2800";
    tmp(57653) := x"2800";
    tmp(57654) := x"2800";
    tmp(57655) := x"2800";
    tmp(57656) := x"2800";
    tmp(57657) := x"2800";
    tmp(57658) := x"2800";
    tmp(57659) := x"2800";
    tmp(57660) := x"2800";
    tmp(57661) := x"2800";
    tmp(57662) := x"2800";
    tmp(57663) := x"2800";
    tmp(57664) := x"2000";
    tmp(57665) := x"2000";
    tmp(57666) := x"2000";
    tmp(57667) := x"2000";
    tmp(57668) := x"2000";
    tmp(57669) := x"1800";
    tmp(57670) := x"1000";
    tmp(57671) := x"1000";
    tmp(57672) := x"0800";
    tmp(57673) := x"0800";
    tmp(57674) := x"0800";
    tmp(57675) := x"0800";
    tmp(57676) := x"0800";
    tmp(57677) := x"1800";
    tmp(57678) := x"1800";
    tmp(57679) := x"1800";
    tmp(57680) := x"2000";
    tmp(57681) := x"2800";
    tmp(57682) := x"2800";
    tmp(57683) := x"2800";
    tmp(57684) := x"2800";
    tmp(57685) := x"2000";
    tmp(57686) := x"2000";
    tmp(57687) := x"2000";
    tmp(57688) := x"2000";
    tmp(57689) := x"2000";
    tmp(57690) := x"1800";
    tmp(57691) := x"1000";
    tmp(57692) := x"1000";
    tmp(57693) := x"1000";
    tmp(57694) := x"1800";
    tmp(57695) := x"2000";
    tmp(57696) := x"1800";
    tmp(57697) := x"1800";
    tmp(57698) := x"2000";
    tmp(57699) := x"2000";
    tmp(57700) := x"2800";
    tmp(57701) := x"2800";
    tmp(57702) := x"3000";
    tmp(57703) := x"3800";
    tmp(57704) := x"4000";
    tmp(57705) := x"4000";
    tmp(57706) := x"4000";
    tmp(57707) := x"3800";
    tmp(57708) := x"3800";
    tmp(57709) := x"3000";
    tmp(57710) := x"3000";
    tmp(57711) := x"3800";
    tmp(57712) := x"4000";
    tmp(57713) := x"4800";
    tmp(57714) := x"5000";
    tmp(57715) := x"5800";
    tmp(57716) := x"6000";
    tmp(57717) := x"5800";
    tmp(57718) := x"5800";
    tmp(57719) := x"5000";
    tmp(57720) := x"5000";
    tmp(57721) := x"5000";
    tmp(57722) := x"5000";
    tmp(57723) := x"5000";
    tmp(57724) := x"5000";
    tmp(57725) := x"5000";
    tmp(57726) := x"5000";
    tmp(57727) := x"5000";
    tmp(57728) := x"5000";
    tmp(57729) := x"5000";
    tmp(57730) := x"5800";
    tmp(57731) := x"5000";
    tmp(57732) := x"4800";
    tmp(57733) := x"4800";
    tmp(57734) := x"5820";
    tmp(57735) := x"5800";
    tmp(57736) := x"5000";
    tmp(57737) := x"7020";
    tmp(57738) := x"6820";
    tmp(57739) := x"6820";
    tmp(57740) := x"7020";
    tmp(57741) := x"6000";
    tmp(57742) := x"5000";
    tmp(57743) := x"5000";
    tmp(57744) := x"5000";
    tmp(57745) := x"5000";
    tmp(57746) := x"5800";
    tmp(57747) := x"5800";
    tmp(57748) := x"6800";
    tmp(57749) := x"6000";
    tmp(57750) := x"8020";
    tmp(57751) := x"7000";
    tmp(57752) := x"7000";
    tmp(57753) := x"7000";
    tmp(57754) := x"7820";
    tmp(57755) := x"7000";
    tmp(57756) := x"7000";
    tmp(57757) := x"8820";
    tmp(57758) := x"8820";
    tmp(57759) := x"7820";
    tmp(57760) := x"6020";
    tmp(57761) := x"6000";
    tmp(57762) := x"5000";
    tmp(57763) := x"3800";
    tmp(57764) := x"4000";
    tmp(57765) := x"4000";
    tmp(57766) := x"5000";
    tmp(57767) := x"6000";
    tmp(57768) := x"6000";
    tmp(57769) := x"6800";
    tmp(57770) := x"8820";
    tmp(57771) := x"a841";
    tmp(57772) := x"b841";
    tmp(57773) := x"c821";
    tmp(57774) := x"b820";
    tmp(57775) := x"b000";
    tmp(57776) := x"b820";
    tmp(57777) := x"a800";
    tmp(57778) := x"9000";
    tmp(57779) := x"c820";
    tmp(57780) := x"c820";
    tmp(57781) := x"a820";
    tmp(57782) := x"c020";
    tmp(57783) := x"d820";
    tmp(57784) := x"e861";
    tmp(57785) := x"6840";
    tmp(57786) := x"1040";
    tmp(57787) := x"0841";
    tmp(57788) := x"0841";
    tmp(57789) := x"0840";
    tmp(57790) := x"0840";
    tmp(57791) := x"0840";
    tmp(57792) := x"0840";
    tmp(57793) := x"0840";
    tmp(57794) := x"0840";
    tmp(57795) := x"0841";
    tmp(57796) := x"0841";
    tmp(57797) := x"0841";
    tmp(57798) := x"0861";
    tmp(57799) := x"0861";
    tmp(57800) := x"1061";
    tmp(57801) := x"1061";
    tmp(57802) := x"1081";
    tmp(57803) := x"1082";
    tmp(57804) := x"1082";
    tmp(57805) := x"1082";
    tmp(57806) := x"10a2";
    tmp(57807) := x"10a2";
    tmp(57808) := x"10a2";
    tmp(57809) := x"10a3";
    tmp(57810) := x"18c3";
    tmp(57811) := x"18c3";
    tmp(57812) := x"18e3";
    tmp(57813) := x"18e3";
    tmp(57814) := x"18e4";
    tmp(57815) := x"18e4";
    tmp(57816) := x"18e4";
    tmp(57817) := x"1904";
    tmp(57818) := x"1904";
    tmp(57819) := x"1903";
    tmp(57820) := x"18e3";
    tmp(57821) := x"18c3";
    tmp(57822) := x"18c3";
    tmp(57823) := x"18c2";
    tmp(57824) := x"10a2";
    tmp(57825) := x"10a2";
    tmp(57826) := x"10a2";
    tmp(57827) := x"1081";
    tmp(57828) := x"1081";
    tmp(57829) := x"1061";
    tmp(57830) := x"0861";
    tmp(57831) := x"0861";
    tmp(57832) := x"0861";
    tmp(57833) := x"0841";
    tmp(57834) := x"0841";
    tmp(57835) := x"0841";
    tmp(57836) := x"0841";
    tmp(57837) := x"0861";
    tmp(57838) := x"0841";
    tmp(57839) := x"0841";
    tmp(57840) := x"0000";
    tmp(57841) := x"0800";
    tmp(57842) := x"0800";
    tmp(57843) := x"0800";
    tmp(57844) := x"0800";
    tmp(57845) := x"0800";
    tmp(57846) := x"0800";
    tmp(57847) := x"0800";
    tmp(57848) := x"0800";
    tmp(57849) := x"0800";
    tmp(57850) := x"0800";
    tmp(57851) := x"1000";
    tmp(57852) := x"1000";
    tmp(57853) := x"1000";
    tmp(57854) := x"0800";
    tmp(57855) := x"0800";
    tmp(57856) := x"0800";
    tmp(57857) := x"1000";
    tmp(57858) := x"1000";
    tmp(57859) := x"1000";
    tmp(57860) := x"1000";
    tmp(57861) := x"1000";
    tmp(57862) := x"1000";
    tmp(57863) := x"1000";
    tmp(57864) := x"1000";
    tmp(57865) := x"1000";
    tmp(57866) := x"1800";
    tmp(57867) := x"1800";
    tmp(57868) := x"1800";
    tmp(57869) := x"1800";
    tmp(57870) := x"1800";
    tmp(57871) := x"1800";
    tmp(57872) := x"1800";
    tmp(57873) := x"1800";
    tmp(57874) := x"2000";
    tmp(57875) := x"2000";
    tmp(57876) := x"2000";
    tmp(57877) := x"2000";
    tmp(57878) := x"2000";
    tmp(57879) := x"2000";
    tmp(57880) := x"2000";
    tmp(57881) := x"2000";
    tmp(57882) := x"2000";
    tmp(57883) := x"2000";
    tmp(57884) := x"2000";
    tmp(57885) := x"2800";
    tmp(57886) := x"2800";
    tmp(57887) := x"2800";
    tmp(57888) := x"2800";
    tmp(57889) := x"2800";
    tmp(57890) := x"2800";
    tmp(57891) := x"2800";
    tmp(57892) := x"2000";
    tmp(57893) := x"2000";
    tmp(57894) := x"2000";
    tmp(57895) := x"2000";
    tmp(57896) := x"2000";
    tmp(57897) := x"2000";
    tmp(57898) := x"2000";
    tmp(57899) := x"2000";
    tmp(57900) := x"2000";
    tmp(57901) := x"2000";
    tmp(57902) := x"2000";
    tmp(57903) := x"2000";
    tmp(57904) := x"2000";
    tmp(57905) := x"2000";
    tmp(57906) := x"1800";
    tmp(57907) := x"1800";
    tmp(57908) := x"2000";
    tmp(57909) := x"2000";
    tmp(57910) := x"2000";
    tmp(57911) := x"1800";
    tmp(57912) := x"1000";
    tmp(57913) := x"1000";
    tmp(57914) := x"1000";
    tmp(57915) := x"1000";
    tmp(57916) := x"1000";
    tmp(57917) := x"1800";
    tmp(57918) := x"2000";
    tmp(57919) := x"2000";
    tmp(57920) := x"2800";
    tmp(57921) := x"2800";
    tmp(57922) := x"2800";
    tmp(57923) := x"2800";
    tmp(57924) := x"2800";
    tmp(57925) := x"2000";
    tmp(57926) := x"1800";
    tmp(57927) := x"2000";
    tmp(57928) := x"1800";
    tmp(57929) := x"2000";
    tmp(57930) := x"1800";
    tmp(57931) := x"1800";
    tmp(57932) := x"1000";
    tmp(57933) := x"1800";
    tmp(57934) := x"2000";
    tmp(57935) := x"2000";
    tmp(57936) := x"2000";
    tmp(57937) := x"2000";
    tmp(57938) := x"2800";
    tmp(57939) := x"3000";
    tmp(57940) := x"3000";
    tmp(57941) := x"2800";
    tmp(57942) := x"2800";
    tmp(57943) := x"3000";
    tmp(57944) := x"3800";
    tmp(57945) := x"3800";
    tmp(57946) := x"4000";
    tmp(57947) := x"4000";
    tmp(57948) := x"3800";
    tmp(57949) := x"3800";
    tmp(57950) := x"3800";
    tmp(57951) := x"3000";
    tmp(57952) := x"3000";
    tmp(57953) := x"3800";
    tmp(57954) := x"4000";
    tmp(57955) := x"5000";
    tmp(57956) := x"5800";
    tmp(57957) := x"5800";
    tmp(57958) := x"5000";
    tmp(57959) := x"5000";
    tmp(57960) := x"5800";
    tmp(57961) := x"5000";
    tmp(57962) := x"5000";
    tmp(57963) := x"5000";
    tmp(57964) := x"5000";
    tmp(57965) := x"5000";
    tmp(57966) := x"5800";
    tmp(57967) := x"5800";
    tmp(57968) := x"5800";
    tmp(57969) := x"5800";
    tmp(57970) := x"6820";
    tmp(57971) := x"6000";
    tmp(57972) := x"5000";
    tmp(57973) := x"5000";
    tmp(57974) := x"5800";
    tmp(57975) := x"5000";
    tmp(57976) := x"5800";
    tmp(57977) := x"8020";
    tmp(57978) := x"6800";
    tmp(57979) := x"7020";
    tmp(57980) := x"7020";
    tmp(57981) := x"5000";
    tmp(57982) := x"5000";
    tmp(57983) := x"5000";
    tmp(57984) := x"5000";
    tmp(57985) := x"4800";
    tmp(57986) := x"5800";
    tmp(57987) := x"5000";
    tmp(57988) := x"6800";
    tmp(57989) := x"6000";
    tmp(57990) := x"7020";
    tmp(57991) := x"7020";
    tmp(57992) := x"8820";
    tmp(57993) := x"7000";
    tmp(57994) := x"7000";
    tmp(57995) := x"7820";
    tmp(57996) := x"8020";
    tmp(57997) := x"8020";
    tmp(57998) := x"9020";
    tmp(57999) := x"8020";
    tmp(58000) := x"7020";
    tmp(58001) := x"6820";
    tmp(58002) := x"6820";
    tmp(58003) := x"3800";
    tmp(58004) := x"4000";
    tmp(58005) := x"5000";
    tmp(58006) := x"5800";
    tmp(58007) := x"6800";
    tmp(58008) := x"6800";
    tmp(58009) := x"7820";
    tmp(58010) := x"9041";
    tmp(58011) := x"a841";
    tmp(58012) := x"d861";
    tmp(58013) := x"f061";
    tmp(58014) := x"d841";
    tmp(58015) := x"d820";
    tmp(58016) := x"d820";
    tmp(58017) := x"d020";
    tmp(58018) := x"9800";
    tmp(58019) := x"f061";
    tmp(58020) := x"b820";
    tmp(58021) := x"a020";
    tmp(58022) := x"b820";
    tmp(58023) := x"d020";
    tmp(58024) := x"d840";
    tmp(58025) := x"5040";
    tmp(58026) := x"1040";
    tmp(58027) := x"0841";
    tmp(58028) := x"0841";
    tmp(58029) := x"0841";
    tmp(58030) := x"0840";
    tmp(58031) := x"0840";
    tmp(58032) := x"0840";
    tmp(58033) := x"0841";
    tmp(58034) := x"0841";
    tmp(58035) := x"0861";
    tmp(58036) := x"0861";
    tmp(58037) := x"1061";
    tmp(58038) := x"1061";
    tmp(58039) := x"1081";
    tmp(58040) := x"1081";
    tmp(58041) := x"1082";
    tmp(58042) := x"10a2";
    tmp(58043) := x"10a2";
    tmp(58044) := x"10a2";
    tmp(58045) := x"10a2";
    tmp(58046) := x"18c3";
    tmp(58047) := x"18c3";
    tmp(58048) := x"18e3";
    tmp(58049) := x"18e3";
    tmp(58050) := x"18e4";
    tmp(58051) := x"18e4";
    tmp(58052) := x"2104";
    tmp(58053) := x"2125";
    tmp(58054) := x"2105";
    tmp(58055) := x"2125";
    tmp(58056) := x"2125";
    tmp(58057) := x"2125";
    tmp(58058) := x"2125";
    tmp(58059) := x"2124";
    tmp(58060) := x"2104";
    tmp(58061) := x"2104";
    tmp(58062) := x"18e4";
    tmp(58063) := x"18e3";
    tmp(58064) := x"18c3";
    tmp(58065) := x"18c3";
    tmp(58066) := x"10c2";
    tmp(58067) := x"10a2";
    tmp(58068) := x"10a2";
    tmp(58069) := x"1081";
    tmp(58070) := x"1081";
    tmp(58071) := x"1061";
    tmp(58072) := x"0861";
    tmp(58073) := x"0861";
    tmp(58074) := x"0861";
    tmp(58075) := x"0861";
    tmp(58076) := x"0861";
    tmp(58077) := x"0861";
    tmp(58078) := x"0861";
    tmp(58079) := x"0861";
    tmp(58080) := x"0000";
    tmp(58081) := x"0800";
    tmp(58082) := x"0800";
    tmp(58083) := x"0800";
    tmp(58084) := x"0800";
    tmp(58085) := x"0800";
    tmp(58086) := x"0800";
    tmp(58087) := x"0800";
    tmp(58088) := x"0800";
    tmp(58089) := x"0800";
    tmp(58090) := x"0800";
    tmp(58091) := x"1000";
    tmp(58092) := x"0800";
    tmp(58093) := x"0800";
    tmp(58094) := x"0800";
    tmp(58095) := x"0800";
    tmp(58096) := x"1000";
    tmp(58097) := x"1000";
    tmp(58098) := x"1000";
    tmp(58099) := x"1000";
    tmp(58100) := x"1000";
    tmp(58101) := x"1000";
    tmp(58102) := x"1000";
    tmp(58103) := x"1000";
    tmp(58104) := x"1000";
    tmp(58105) := x"1000";
    tmp(58106) := x"1800";
    tmp(58107) := x"1800";
    tmp(58108) := x"1800";
    tmp(58109) := x"1800";
    tmp(58110) := x"1800";
    tmp(58111) := x"1800";
    tmp(58112) := x"2000";
    tmp(58113) := x"2000";
    tmp(58114) := x"2000";
    tmp(58115) := x"2800";
    tmp(58116) := x"2000";
    tmp(58117) := x"2000";
    tmp(58118) := x"2000";
    tmp(58119) := x"2000";
    tmp(58120) := x"2000";
    tmp(58121) := x"2000";
    tmp(58122) := x"2000";
    tmp(58123) := x"2000";
    tmp(58124) := x"2000";
    tmp(58125) := x"2800";
    tmp(58126) := x"2800";
    tmp(58127) := x"2800";
    tmp(58128) := x"2800";
    tmp(58129) := x"2800";
    tmp(58130) := x"2800";
    tmp(58131) := x"2800";
    tmp(58132) := x"2000";
    tmp(58133) := x"2000";
    tmp(58134) := x"1800";
    tmp(58135) := x"1800";
    tmp(58136) := x"2000";
    tmp(58137) := x"2000";
    tmp(58138) := x"1800";
    tmp(58139) := x"1800";
    tmp(58140) := x"1800";
    tmp(58141) := x"2000";
    tmp(58142) := x"2000";
    tmp(58143) := x"2800";
    tmp(58144) := x"2800";
    tmp(58145) := x"2000";
    tmp(58146) := x"1800";
    tmp(58147) := x"1800";
    tmp(58148) := x"1800";
    tmp(58149) := x"1800";
    tmp(58150) := x"2000";
    tmp(58151) := x"2000";
    tmp(58152) := x"2000";
    tmp(58153) := x"1800";
    tmp(58154) := x"1800";
    tmp(58155) := x"1800";
    tmp(58156) := x"1800";
    tmp(58157) := x"1800";
    tmp(58158) := x"2800";
    tmp(58159) := x"2800";
    tmp(58160) := x"2800";
    tmp(58161) := x"3000";
    tmp(58162) := x"2800";
    tmp(58163) := x"2800";
    tmp(58164) := x"2800";
    tmp(58165) := x"2000";
    tmp(58166) := x"1800";
    tmp(58167) := x"1800";
    tmp(58168) := x"1800";
    tmp(58169) := x"1800";
    tmp(58170) := x"2000";
    tmp(58171) := x"2000";
    tmp(58172) := x"1800";
    tmp(58173) := x"1800";
    tmp(58174) := x"2000";
    tmp(58175) := x"2000";
    tmp(58176) := x"2000";
    tmp(58177) := x"2800";
    tmp(58178) := x"2800";
    tmp(58179) := x"3000";
    tmp(58180) := x"2800";
    tmp(58181) := x"2800";
    tmp(58182) := x"2800";
    tmp(58183) := x"3000";
    tmp(58184) := x"3800";
    tmp(58185) := x"4000";
    tmp(58186) := x"4000";
    tmp(58187) := x"4000";
    tmp(58188) := x"4000";
    tmp(58189) := x"3800";
    tmp(58190) := x"3800";
    tmp(58191) := x"3000";
    tmp(58192) := x"2800";
    tmp(58193) := x"2800";
    tmp(58194) := x"3000";
    tmp(58195) := x"4000";
    tmp(58196) := x"4000";
    tmp(58197) := x"4800";
    tmp(58198) := x"5000";
    tmp(58199) := x"5800";
    tmp(58200) := x"5000";
    tmp(58201) := x"5000";
    tmp(58202) := x"5000";
    tmp(58203) := x"5000";
    tmp(58204) := x"5000";
    tmp(58205) := x"5000";
    tmp(58206) := x"5800";
    tmp(58207) := x"5800";
    tmp(58208) := x"5800";
    tmp(58209) := x"6000";
    tmp(58210) := x"6800";
    tmp(58211) := x"6000";
    tmp(58212) := x"5000";
    tmp(58213) := x"5000";
    tmp(58214) := x"5000";
    tmp(58215) := x"5000";
    tmp(58216) := x"6000";
    tmp(58217) := x"7020";
    tmp(58218) := x"6800";
    tmp(58219) := x"7020";
    tmp(58220) := x"7020";
    tmp(58221) := x"5000";
    tmp(58222) := x"5000";
    tmp(58223) := x"5000";
    tmp(58224) := x"5800";
    tmp(58225) := x"5000";
    tmp(58226) := x"5800";
    tmp(58227) := x"5000";
    tmp(58228) := x"6820";
    tmp(58229) := x"6820";
    tmp(58230) := x"6820";
    tmp(58231) := x"7820";
    tmp(58232) := x"8820";
    tmp(58233) := x"7000";
    tmp(58234) := x"7000";
    tmp(58235) := x"7820";
    tmp(58236) := x"8820";
    tmp(58237) := x"8020";
    tmp(58238) := x"8820";
    tmp(58239) := x"8020";
    tmp(58240) := x"7820";
    tmp(58241) := x"7020";
    tmp(58242) := x"7020";
    tmp(58243) := x"4000";
    tmp(58244) := x"4000";
    tmp(58245) := x"5000";
    tmp(58246) := x"6000";
    tmp(58247) := x"7000";
    tmp(58248) := x"6800";
    tmp(58249) := x"9021";
    tmp(58250) := x"a061";
    tmp(58251) := x"a861";
    tmp(58252) := x"c861";
    tmp(58253) := x"d041";
    tmp(58254) := x"d841";
    tmp(58255) := x"f881";
    tmp(58256) := x"e820";
    tmp(58257) := x"e020";
    tmp(58258) := x"a000";
    tmp(58259) := x"f861";
    tmp(58260) := x"b020";
    tmp(58261) := x"a800";
    tmp(58262) := x"c020";
    tmp(58263) := x"c820";
    tmp(58264) := x"c840";
    tmp(58265) := x"4061";
    tmp(58266) := x"0840";
    tmp(58267) := x"0841";
    tmp(58268) := x"0841";
    tmp(58269) := x"0841";
    tmp(58270) := x"0841";
    tmp(58271) := x"0841";
    tmp(58272) := x"0841";
    tmp(58273) := x"0861";
    tmp(58274) := x"1061";
    tmp(58275) := x"1061";
    tmp(58276) := x"1061";
    tmp(58277) := x"1081";
    tmp(58278) := x"1082";
    tmp(58279) := x"1082";
    tmp(58280) := x"10a2";
    tmp(58281) := x"10a2";
    tmp(58282) := x"18a2";
    tmp(58283) := x"18a3";
    tmp(58284) := x"18c3";
    tmp(58285) := x"18c3";
    tmp(58286) := x"18e4";
    tmp(58287) := x"2104";
    tmp(58288) := x"2104";
    tmp(58289) := x"2104";
    tmp(58290) := x"2125";
    tmp(58291) := x"2125";
    tmp(58292) := x"2945";
    tmp(58293) := x"2945";
    tmp(58294) := x"2946";
    tmp(58295) := x"2946";
    tmp(58296) := x"2946";
    tmp(58297) := x"2946";
    tmp(58298) := x"2946";
    tmp(58299) := x"2946";
    tmp(58300) := x"2946";
    tmp(58301) := x"2125";
    tmp(58302) := x"2124";
    tmp(58303) := x"2104";
    tmp(58304) := x"2104";
    tmp(58305) := x"18e3";
    tmp(58306) := x"18e3";
    tmp(58307) := x"18c3";
    tmp(58308) := x"10a2";
    tmp(58309) := x"10a2";
    tmp(58310) := x"10a1";
    tmp(58311) := x"1081";
    tmp(58312) := x"1081";
    tmp(58313) := x"0861";
    tmp(58314) := x"0861";
    tmp(58315) := x"0861";
    tmp(58316) := x"0861";
    tmp(58317) := x"0861";
    tmp(58318) := x"0861";
    tmp(58319) := x"0861";
    tmp(58320) := x"0000";
    tmp(58321) := x"1000";
    tmp(58322) := x"1000";
    tmp(58323) := x"0800";
    tmp(58324) := x"0800";
    tmp(58325) := x"0800";
    tmp(58326) := x"0800";
    tmp(58327) := x"0800";
    tmp(58328) := x"0800";
    tmp(58329) := x"0800";
    tmp(58330) := x"0800";
    tmp(58331) := x"0800";
    tmp(58332) := x"0800";
    tmp(58333) := x"0800";
    tmp(58334) := x"0800";
    tmp(58335) := x"0800";
    tmp(58336) := x"1000";
    tmp(58337) := x"1000";
    tmp(58338) := x"1000";
    tmp(58339) := x"1000";
    tmp(58340) := x"1000";
    tmp(58341) := x"1000";
    tmp(58342) := x"1000";
    tmp(58343) := x"1000";
    tmp(58344) := x"1000";
    tmp(58345) := x"1000";
    tmp(58346) := x"1800";
    tmp(58347) := x"1800";
    tmp(58348) := x"1800";
    tmp(58349) := x"1800";
    tmp(58350) := x"1800";
    tmp(58351) := x"2000";
    tmp(58352) := x"2000";
    tmp(58353) := x"2000";
    tmp(58354) := x"2000";
    tmp(58355) := x"2000";
    tmp(58356) := x"2000";
    tmp(58357) := x"2000";
    tmp(58358) := x"2000";
    tmp(58359) := x"2000";
    tmp(58360) := x"2000";
    tmp(58361) := x"2000";
    tmp(58362) := x"2000";
    tmp(58363) := x"2000";
    tmp(58364) := x"2800";
    tmp(58365) := x"2800";
    tmp(58366) := x"2800";
    tmp(58367) := x"2800";
    tmp(58368) := x"2800";
    tmp(58369) := x"2800";
    tmp(58370) := x"2800";
    tmp(58371) := x"2000";
    tmp(58372) := x"2000";
    tmp(58373) := x"2000";
    tmp(58374) := x"1800";
    tmp(58375) := x"1800";
    tmp(58376) := x"2000";
    tmp(58377) := x"2000";
    tmp(58378) := x"2000";
    tmp(58379) := x"2000";
    tmp(58380) := x"2000";
    tmp(58381) := x"2000";
    tmp(58382) := x"2800";
    tmp(58383) := x"2800";
    tmp(58384) := x"2800";
    tmp(58385) := x"2800";
    tmp(58386) := x"2800";
    tmp(58387) := x"2000";
    tmp(58388) := x"2000";
    tmp(58389) := x"1800";
    tmp(58390) := x"1000";
    tmp(58391) := x"1000";
    tmp(58392) := x"1000";
    tmp(58393) := x"1000";
    tmp(58394) := x"1000";
    tmp(58395) := x"1800";
    tmp(58396) := x"1800";
    tmp(58397) := x"1800";
    tmp(58398) := x"2000";
    tmp(58399) := x"2000";
    tmp(58400) := x"2800";
    tmp(58401) := x"2800";
    tmp(58402) := x"2800";
    tmp(58403) := x"2800";
    tmp(58404) := x"2800";
    tmp(58405) := x"2000";
    tmp(58406) := x"1800";
    tmp(58407) := x"1800";
    tmp(58408) := x"2000";
    tmp(58409) := x"2000";
    tmp(58410) := x"2000";
    tmp(58411) := x"2000";
    tmp(58412) := x"2000";
    tmp(58413) := x"1800";
    tmp(58414) := x"1800";
    tmp(58415) := x"2000";
    tmp(58416) := x"2800";
    tmp(58417) := x"3000";
    tmp(58418) := x"3000";
    tmp(58419) := x"3000";
    tmp(58420) := x"2800";
    tmp(58421) := x"2000";
    tmp(58422) := x"2800";
    tmp(58423) := x"3000";
    tmp(58424) := x"3800";
    tmp(58425) := x"4000";
    tmp(58426) := x"4000";
    tmp(58427) := x"4800";
    tmp(58428) := x"4800";
    tmp(58429) := x"4000";
    tmp(58430) := x"4000";
    tmp(58431) := x"3800";
    tmp(58432) := x"3000";
    tmp(58433) := x"3000";
    tmp(58434) := x"3800";
    tmp(58435) := x"3800";
    tmp(58436) := x"4000";
    tmp(58437) := x"4800";
    tmp(58438) := x"5000";
    tmp(58439) := x"4000";
    tmp(58440) := x"3800";
    tmp(58441) := x"5000";
    tmp(58442) := x"5000";
    tmp(58443) := x"5000";
    tmp(58444) := x"4800";
    tmp(58445) := x"4800";
    tmp(58446) := x"5000";
    tmp(58447) := x"5000";
    tmp(58448) := x"5800";
    tmp(58449) := x"5800";
    tmp(58450) := x"6000";
    tmp(58451) := x"6000";
    tmp(58452) := x"5800";
    tmp(58453) := x"5000";
    tmp(58454) := x"5000";
    tmp(58455) := x"5000";
    tmp(58456) := x"6800";
    tmp(58457) := x"6800";
    tmp(58458) := x"6000";
    tmp(58459) := x"7020";
    tmp(58460) := x"6800";
    tmp(58461) := x"5000";
    tmp(58462) := x"5000";
    tmp(58463) := x"5000";
    tmp(58464) := x"5800";
    tmp(58465) := x"5800";
    tmp(58466) := x"5800";
    tmp(58467) := x"5800";
    tmp(58468) := x"6020";
    tmp(58469) := x"7020";
    tmp(58470) := x"6020";
    tmp(58471) := x"7820";
    tmp(58472) := x"7820";
    tmp(58473) := x"8020";
    tmp(58474) := x"7820";
    tmp(58475) := x"7020";
    tmp(58476) := x"8020";
    tmp(58477) := x"8820";
    tmp(58478) := x"7820";
    tmp(58479) := x"8020";
    tmp(58480) := x"8820";
    tmp(58481) := x"7820";
    tmp(58482) := x"7820";
    tmp(58483) := x"5800";
    tmp(58484) := x"4000";
    tmp(58485) := x"5800";
    tmp(58486) := x"6800";
    tmp(58487) := x"8820";
    tmp(58488) := x"9020";
    tmp(58489) := x"a841";
    tmp(58490) := x"c082";
    tmp(58491) := x"b862";
    tmp(58492) := x"b041";
    tmp(58493) := x"a021";
    tmp(58494) := x"d861";
    tmp(58495) := x"e861";
    tmp(58496) := x"e020";
    tmp(58497) := x"d820";
    tmp(58498) := x"a820";
    tmp(58499) := x"f860";
    tmp(58500) := x"c020";
    tmp(58501) := x"a820";
    tmp(58502) := x"c020";
    tmp(58503) := x"b020";
    tmp(58504) := x"a840";
    tmp(58505) := x"3061";
    tmp(58506) := x"0840";
    tmp(58507) := x"0841";
    tmp(58508) := x"0841";
    tmp(58509) := x"0841";
    tmp(58510) := x"0841";
    tmp(58511) := x"0841";
    tmp(58512) := x"0861";
    tmp(58513) := x"1061";
    tmp(58514) := x"1061";
    tmp(58515) := x"1081";
    tmp(58516) := x"1081";
    tmp(58517) := x"10a2";
    tmp(58518) := x"10a2";
    tmp(58519) := x"18a2";
    tmp(58520) := x"18c2";
    tmp(58521) := x"18c3";
    tmp(58522) := x"18c3";
    tmp(58523) := x"18e3";
    tmp(58524) := x"18e4";
    tmp(58525) := x"2104";
    tmp(58526) := x"2104";
    tmp(58527) := x"2125";
    tmp(58528) := x"2125";
    tmp(58529) := x"2125";
    tmp(58530) := x"2946";
    tmp(58531) := x"2946";
    tmp(58532) := x"2946";
    tmp(58533) := x"2966";
    tmp(58534) := x"2966";
    tmp(58535) := x"2967";
    tmp(58536) := x"2967";
    tmp(58537) := x"2967";
    tmp(58538) := x"2967";
    tmp(58539) := x"2987";
    tmp(58540) := x"2967";
    tmp(58541) := x"2966";
    tmp(58542) := x"2945";
    tmp(58543) := x"2945";
    tmp(58544) := x"2125";
    tmp(58545) := x"2104";
    tmp(58546) := x"2104";
    tmp(58547) := x"18e3";
    tmp(58548) := x"18c3";
    tmp(58549) := x"18c2";
    tmp(58550) := x"10c2";
    tmp(58551) := x"10a2";
    tmp(58552) := x"1081";
    tmp(58553) := x"1081";
    tmp(58554) := x"1081";
    tmp(58555) := x"0861";
    tmp(58556) := x"0861";
    tmp(58557) := x"0861";
    tmp(58558) := x"0861";
    tmp(58559) := x"0861";
    tmp(58560) := x"0000";
    tmp(58561) := x"1000";
    tmp(58562) := x"1000";
    tmp(58563) := x"0800";
    tmp(58564) := x"0800";
    tmp(58565) := x"0800";
    tmp(58566) := x"0800";
    tmp(58567) := x"0800";
    tmp(58568) := x"0800";
    tmp(58569) := x"0800";
    tmp(58570) := x"0800";
    tmp(58571) := x"0800";
    tmp(58572) := x"0800";
    tmp(58573) := x"0800";
    tmp(58574) := x"1000";
    tmp(58575) := x"1000";
    tmp(58576) := x"1000";
    tmp(58577) := x"1000";
    tmp(58578) := x"1000";
    tmp(58579) := x"1000";
    tmp(58580) := x"1000";
    tmp(58581) := x"1800";
    tmp(58582) := x"1000";
    tmp(58583) := x"1000";
    tmp(58584) := x"1000";
    tmp(58585) := x"1000";
    tmp(58586) := x"1800";
    tmp(58587) := x"1800";
    tmp(58588) := x"1800";
    tmp(58589) := x"1800";
    tmp(58590) := x"1800";
    tmp(58591) := x"2000";
    tmp(58592) := x"2000";
    tmp(58593) := x"2000";
    tmp(58594) := x"2000";
    tmp(58595) := x"2000";
    tmp(58596) := x"2000";
    tmp(58597) := x"1800";
    tmp(58598) := x"2000";
    tmp(58599) := x"2000";
    tmp(58600) := x"2000";
    tmp(58601) := x"2000";
    tmp(58602) := x"2800";
    tmp(58603) := x"2000";
    tmp(58604) := x"2800";
    tmp(58605) := x"2800";
    tmp(58606) := x"2800";
    tmp(58607) := x"2800";
    tmp(58608) := x"2800";
    tmp(58609) := x"2800";
    tmp(58610) := x"2000";
    tmp(58611) := x"2000";
    tmp(58612) := x"2000";
    tmp(58613) := x"2000";
    tmp(58614) := x"2000";
    tmp(58615) := x"2800";
    tmp(58616) := x"2800";
    tmp(58617) := x"2000";
    tmp(58618) := x"2800";
    tmp(58619) := x"2800";
    tmp(58620) := x"2800";
    tmp(58621) := x"2800";
    tmp(58622) := x"2800";
    tmp(58623) := x"2800";
    tmp(58624) := x"2800";
    tmp(58625) := x"2800";
    tmp(58626) := x"2800";
    tmp(58627) := x"2800";
    tmp(58628) := x"2000";
    tmp(58629) := x"2000";
    tmp(58630) := x"1800";
    tmp(58631) := x"0800";
    tmp(58632) := x"0800";
    tmp(58633) := x"0800";
    tmp(58634) := x"0800";
    tmp(58635) := x"1000";
    tmp(58636) := x"1000";
    tmp(58637) := x"1000";
    tmp(58638) := x"1800";
    tmp(58639) := x"2000";
    tmp(58640) := x"2000";
    tmp(58641) := x"2800";
    tmp(58642) := x"2800";
    tmp(58643) := x"2800";
    tmp(58644) := x"2800";
    tmp(58645) := x"2000";
    tmp(58646) := x"1800";
    tmp(58647) := x"1800";
    tmp(58648) := x"1800";
    tmp(58649) := x"1800";
    tmp(58650) := x"1000";
    tmp(58651) := x"1800";
    tmp(58652) := x"2000";
    tmp(58653) := x"2000";
    tmp(58654) := x"1800";
    tmp(58655) := x"2000";
    tmp(58656) := x"2800";
    tmp(58657) := x"3000";
    tmp(58658) := x"3000";
    tmp(58659) := x"3000";
    tmp(58660) := x"2800";
    tmp(58661) := x"2800";
    tmp(58662) := x"2800";
    tmp(58663) := x"3000";
    tmp(58664) := x"3800";
    tmp(58665) := x"4000";
    tmp(58666) := x"4000";
    tmp(58667) := x"4000";
    tmp(58668) := x"4000";
    tmp(58669) := x"4800";
    tmp(58670) := x"5000";
    tmp(58671) := x"5000";
    tmp(58672) := x"4800";
    tmp(58673) := x"4000";
    tmp(58674) := x"3800";
    tmp(58675) := x"3000";
    tmp(58676) := x"3000";
    tmp(58677) := x"3800";
    tmp(58678) := x"3000";
    tmp(58679) := x"2800";
    tmp(58680) := x"4000";
    tmp(58681) := x"5000";
    tmp(58682) := x"5000";
    tmp(58683) := x"4800";
    tmp(58684) := x"4800";
    tmp(58685) := x"5000";
    tmp(58686) := x"5800";
    tmp(58687) := x"5800";
    tmp(58688) := x"5800";
    tmp(58689) := x"5800";
    tmp(58690) := x"6800";
    tmp(58691) := x"6800";
    tmp(58692) := x"6000";
    tmp(58693) := x"5800";
    tmp(58694) := x"5000";
    tmp(58695) := x"5800";
    tmp(58696) := x"6820";
    tmp(58697) := x"6000";
    tmp(58698) := x"6000";
    tmp(58699) := x"7000";
    tmp(58700) := x"6000";
    tmp(58701) := x"5000";
    tmp(58702) := x"5000";
    tmp(58703) := x"5000";
    tmp(58704) := x"5800";
    tmp(58705) := x"5800";
    tmp(58706) := x"5800";
    tmp(58707) := x"6000";
    tmp(58708) := x"5800";
    tmp(58709) := x"7820";
    tmp(58710) := x"6020";
    tmp(58711) := x"6820";
    tmp(58712) := x"7820";
    tmp(58713) := x"8820";
    tmp(58714) := x"7820";
    tmp(58715) := x"7820";
    tmp(58716) := x"7820";
    tmp(58717) := x"8820";
    tmp(58718) := x"8020";
    tmp(58719) := x"8820";
    tmp(58720) := x"8020";
    tmp(58721) := x"9020";
    tmp(58722) := x"7820";
    tmp(58723) := x"6800";
    tmp(58724) := x"4800";
    tmp(58725) := x"5800";
    tmp(58726) := x"7000";
    tmp(58727) := x"a020";
    tmp(58728) := x"b841";
    tmp(58729) := x"c881";
    tmp(58730) := x"d0a2";
    tmp(58731) := x"e904";
    tmp(58732) := x"d0c3";
    tmp(58733) := x"b062";
    tmp(58734) := x"d8a2";
    tmp(58735) := x"d841";
    tmp(58736) := x"e820";
    tmp(58737) := x"c820";
    tmp(58738) := x"c020";
    tmp(58739) := x"f040";
    tmp(58740) := x"c820";
    tmp(58741) := x"b820";
    tmp(58742) := x"c820";
    tmp(58743) := x"a020";
    tmp(58744) := x"9041";
    tmp(58745) := x"2061";
    tmp(58746) := x"0840";
    tmp(58747) := x"0841";
    tmp(58748) := x"0841";
    tmp(58749) := x"0841";
    tmp(58750) := x"0861";
    tmp(58751) := x"1061";
    tmp(58752) := x"1061";
    tmp(58753) := x"1061";
    tmp(58754) := x"1081";
    tmp(58755) := x"10a2";
    tmp(58756) := x"10a2";
    tmp(58757) := x"10a2";
    tmp(58758) := x"18c3";
    tmp(58759) := x"18c3";
    tmp(58760) := x"18c3";
    tmp(58761) := x"18e3";
    tmp(58762) := x"20e4";
    tmp(58763) := x"2104";
    tmp(58764) := x"2104";
    tmp(58765) := x"2125";
    tmp(58766) := x"2125";
    tmp(58767) := x"2945";
    tmp(58768) := x"2946";
    tmp(58769) := x"2946";
    tmp(58770) := x"2966";
    tmp(58771) := x"2966";
    tmp(58772) := x"2987";
    tmp(58773) := x"2987";
    tmp(58774) := x"2967";
    tmp(58775) := x"3187";
    tmp(58776) := x"3187";
    tmp(58777) := x"3187";
    tmp(58778) := x"31a7";
    tmp(58779) := x"31a7";
    tmp(58780) := x"3187";
    tmp(58781) := x"31a7";
    tmp(58782) := x"3187";
    tmp(58783) := x"2966";
    tmp(58784) := x"2965";
    tmp(58785) := x"2945";
    tmp(58786) := x"2125";
    tmp(58787) := x"2104";
    tmp(58788) := x"1903";
    tmp(58789) := x"18e3";
    tmp(58790) := x"18c3";
    tmp(58791) := x"10a2";
    tmp(58792) := x"10a2";
    tmp(58793) := x"1081";
    tmp(58794) := x"1081";
    tmp(58795) := x"1061";
    tmp(58796) := x"0861";
    tmp(58797) := x"0861";
    tmp(58798) := x"0861";
    tmp(58799) := x"0861";
    tmp(58800) := x"0000";
    tmp(58801) := x"0800";
    tmp(58802) := x"0800";
    tmp(58803) := x"0800";
    tmp(58804) := x"0800";
    tmp(58805) := x"0800";
    tmp(58806) := x"0800";
    tmp(58807) := x"0800";
    tmp(58808) := x"0800";
    tmp(58809) := x"0800";
    tmp(58810) := x"0800";
    tmp(58811) := x"0800";
    tmp(58812) := x"1000";
    tmp(58813) := x"1000";
    tmp(58814) := x"1000";
    tmp(58815) := x"1000";
    tmp(58816) := x"1000";
    tmp(58817) := x"1000";
    tmp(58818) := x"1000";
    tmp(58819) := x"1000";
    tmp(58820) := x"1000";
    tmp(58821) := x"1000";
    tmp(58822) := x"1000";
    tmp(58823) := x"1000";
    tmp(58824) := x"1000";
    tmp(58825) := x"1000";
    tmp(58826) := x"1000";
    tmp(58827) := x"1800";
    tmp(58828) := x"1800";
    tmp(58829) := x"1800";
    tmp(58830) := x"2000";
    tmp(58831) := x"2000";
    tmp(58832) := x"2000";
    tmp(58833) := x"2000";
    tmp(58834) := x"2000";
    tmp(58835) := x"2000";
    tmp(58836) := x"2000";
    tmp(58837) := x"1800";
    tmp(58838) := x"1800";
    tmp(58839) := x"2000";
    tmp(58840) := x"2000";
    tmp(58841) := x"2000";
    tmp(58842) := x"2800";
    tmp(58843) := x"2000";
    tmp(58844) := x"2000";
    tmp(58845) := x"2800";
    tmp(58846) := x"2800";
    tmp(58847) := x"2800";
    tmp(58848) := x"2800";
    tmp(58849) := x"2800";
    tmp(58850) := x"2800";
    tmp(58851) := x"3000";
    tmp(58852) := x"3000";
    tmp(58853) := x"3000";
    tmp(58854) := x"2800";
    tmp(58855) := x"2800";
    tmp(58856) := x"2800";
    tmp(58857) := x"2800";
    tmp(58858) := x"2800";
    tmp(58859) := x"2800";
    tmp(58860) := x"2800";
    tmp(58861) := x"2800";
    tmp(58862) := x"2800";
    tmp(58863) := x"2800";
    tmp(58864) := x"2800";
    tmp(58865) := x"2800";
    tmp(58866) := x"2800";
    tmp(58867) := x"2800";
    tmp(58868) := x"2000";
    tmp(58869) := x"2000";
    tmp(58870) := x"1800";
    tmp(58871) := x"1000";
    tmp(58872) := x"1000";
    tmp(58873) := x"0800";
    tmp(58874) := x"0800";
    tmp(58875) := x"1000";
    tmp(58876) := x"1000";
    tmp(58877) := x"1800";
    tmp(58878) := x"1800";
    tmp(58879) := x"2000";
    tmp(58880) := x"2000";
    tmp(58881) := x"2000";
    tmp(58882) := x"2000";
    tmp(58883) := x"2000";
    tmp(58884) := x"2000";
    tmp(58885) := x"2000";
    tmp(58886) := x"1800";
    tmp(58887) := x"1000";
    tmp(58888) := x"1000";
    tmp(58889) := x"1000";
    tmp(58890) := x"1800";
    tmp(58891) := x"2000";
    tmp(58892) := x"2000";
    tmp(58893) := x"2000";
    tmp(58894) := x"2000";
    tmp(58895) := x"2000";
    tmp(58896) := x"2800";
    tmp(58897) := x"2800";
    tmp(58898) := x"3000";
    tmp(58899) := x"3000";
    tmp(58900) := x"2800";
    tmp(58901) := x"3000";
    tmp(58902) := x"3800";
    tmp(58903) := x"3800";
    tmp(58904) := x"4000";
    tmp(58905) := x"4000";
    tmp(58906) := x"4000";
    tmp(58907) := x"4800";
    tmp(58908) := x"4800";
    tmp(58909) := x"4800";
    tmp(58910) := x"5000";
    tmp(58911) := x"5000";
    tmp(58912) := x"4800";
    tmp(58913) := x"4000";
    tmp(58914) := x"4000";
    tmp(58915) := x"3800";
    tmp(58916) := x"3000";
    tmp(58917) := x"2800";
    tmp(58918) := x"2800";
    tmp(58919) := x"4000";
    tmp(58920) := x"4800";
    tmp(58921) := x"4800";
    tmp(58922) := x"4800";
    tmp(58923) := x"4800";
    tmp(58924) := x"4800";
    tmp(58925) := x"5800";
    tmp(58926) := x"6000";
    tmp(58927) := x"5800";
    tmp(58928) := x"5800";
    tmp(58929) := x"6000";
    tmp(58930) := x"6800";
    tmp(58931) := x"6000";
    tmp(58932) := x"6000";
    tmp(58933) := x"6000";
    tmp(58934) := x"5800";
    tmp(58935) := x"6000";
    tmp(58936) := x"7020";
    tmp(58937) := x"5800";
    tmp(58938) := x"6000";
    tmp(58939) := x"7000";
    tmp(58940) := x"5800";
    tmp(58941) := x"5000";
    tmp(58942) := x"5800";
    tmp(58943) := x"5000";
    tmp(58944) := x"5800";
    tmp(58945) := x"5800";
    tmp(58946) := x"5800";
    tmp(58947) := x"5800";
    tmp(58948) := x"6020";
    tmp(58949) := x"8020";
    tmp(58950) := x"6820";
    tmp(58951) := x"6820";
    tmp(58952) := x"7020";
    tmp(58953) := x"7820";
    tmp(58954) := x"7820";
    tmp(58955) := x"7820";
    tmp(58956) := x"7020";
    tmp(58957) := x"8820";
    tmp(58958) := x"8820";
    tmp(58959) := x"8820";
    tmp(58960) := x"7820";
    tmp(58961) := x"a840";
    tmp(58962) := x"8020";
    tmp(58963) := x"7000";
    tmp(58964) := x"5000";
    tmp(58965) := x"6000";
    tmp(58966) := x"7800";
    tmp(58967) := x"a020";
    tmp(58968) := x"c041";
    tmp(58969) := x"e081";
    tmp(58970) := x"f0e3";
    tmp(58971) := x"f9a7";
    tmp(58972) := x"f1c8";
    tmp(58973) := x"e125";
    tmp(58974) := x"e8c3";
    tmp(58975) := x"e861";
    tmp(58976) := x"f841";
    tmp(58977) := x"b020";
    tmp(58978) := x"d020";
    tmp(58979) := x"f040";
    tmp(58980) := x"d020";
    tmp(58981) := x"c820";
    tmp(58982) := x"b020";
    tmp(58983) := x"a820";
    tmp(58984) := x"6061";
    tmp(58985) := x"1040";
    tmp(58986) := x"0841";
    tmp(58987) := x"0841";
    tmp(58988) := x"0841";
    tmp(58989) := x"0861";
    tmp(58990) := x"1061";
    tmp(58991) := x"1061";
    tmp(58992) := x"1081";
    tmp(58993) := x"1081";
    tmp(58994) := x"10a2";
    tmp(58995) := x"10a2";
    tmp(58996) := x"18a2";
    tmp(58997) := x"18c3";
    tmp(58998) := x"18e3";
    tmp(58999) := x"18e3";
    tmp(59000) := x"18e4";
    tmp(59001) := x"20e4";
    tmp(59002) := x"2104";
    tmp(59003) := x"2124";
    tmp(59004) := x"2925";
    tmp(59005) := x"2945";
    tmp(59006) := x"2946";
    tmp(59007) := x"2966";
    tmp(59008) := x"2967";
    tmp(59009) := x"3187";
    tmp(59010) := x"3187";
    tmp(59011) := x"3187";
    tmp(59012) := x"31a7";
    tmp(59013) := x"31a8";
    tmp(59014) := x"31a8";
    tmp(59015) := x"31a8";
    tmp(59016) := x"39c8";
    tmp(59017) := x"31c8";
    tmp(59018) := x"31a8";
    tmp(59019) := x"31a8";
    tmp(59020) := x"39c8";
    tmp(59021) := x"39c8";
    tmp(59022) := x"31c8";
    tmp(59023) := x"31a7";
    tmp(59024) := x"3186";
    tmp(59025) := x"2966";
    tmp(59026) := x"2945";
    tmp(59027) := x"2945";
    tmp(59028) := x"2124";
    tmp(59029) := x"1903";
    tmp(59030) := x"18e3";
    tmp(59031) := x"10c2";
    tmp(59032) := x"10a2";
    tmp(59033) := x"1081";
    tmp(59034) := x"1081";
    tmp(59035) := x"0861";
    tmp(59036) := x"0861";
    tmp(59037) := x"0861";
    tmp(59038) := x"0861";
    tmp(59039) := x"0861";
    tmp(59040) := x"0000";
    tmp(59041) := x"0800";
    tmp(59042) := x"0800";
    tmp(59043) := x"0800";
    tmp(59044) := x"0800";
    tmp(59045) := x"0800";
    tmp(59046) := x"0800";
    tmp(59047) := x"0800";
    tmp(59048) := x"0800";
    tmp(59049) := x"0800";
    tmp(59050) := x"0800";
    tmp(59051) := x"1000";
    tmp(59052) := x"1000";
    tmp(59053) := x"1000";
    tmp(59054) := x"1000";
    tmp(59055) := x"1000";
    tmp(59056) := x"1000";
    tmp(59057) := x"1000";
    tmp(59058) := x"1000";
    tmp(59059) := x"1000";
    tmp(59060) := x"1000";
    tmp(59061) := x"1800";
    tmp(59062) := x"1000";
    tmp(59063) := x"1000";
    tmp(59064) := x"1000";
    tmp(59065) := x"1000";
    tmp(59066) := x"1800";
    tmp(59067) := x"1800";
    tmp(59068) := x"1800";
    tmp(59069) := x"2000";
    tmp(59070) := x"2000";
    tmp(59071) := x"2000";
    tmp(59072) := x"2000";
    tmp(59073) := x"2000";
    tmp(59074) := x"2000";
    tmp(59075) := x"2000";
    tmp(59076) := x"2000";
    tmp(59077) := x"2000";
    tmp(59078) := x"2000";
    tmp(59079) := x"2000";
    tmp(59080) := x"2000";
    tmp(59081) := x"2800";
    tmp(59082) := x"2800";
    tmp(59083) := x"2000";
    tmp(59084) := x"2000";
    tmp(59085) := x"2800";
    tmp(59086) := x"2800";
    tmp(59087) := x"2800";
    tmp(59088) := x"2800";
    tmp(59089) := x"2800";
    tmp(59090) := x"2800";
    tmp(59091) := x"3000";
    tmp(59092) := x"3000";
    tmp(59093) := x"3000";
    tmp(59094) := x"2800";
    tmp(59095) := x"2800";
    tmp(59096) := x"2800";
    tmp(59097) := x"2800";
    tmp(59098) := x"2800";
    tmp(59099) := x"2800";
    tmp(59100) := x"2800";
    tmp(59101) := x"2800";
    tmp(59102) := x"2800";
    tmp(59103) := x"2800";
    tmp(59104) := x"2800";
    tmp(59105) := x"2800";
    tmp(59106) := x"2800";
    tmp(59107) := x"2000";
    tmp(59108) := x"2000";
    tmp(59109) := x"2000";
    tmp(59110) := x"1800";
    tmp(59111) := x"1800";
    tmp(59112) := x"1000";
    tmp(59113) := x"1000";
    tmp(59114) := x"1000";
    tmp(59115) := x"1000";
    tmp(59116) := x"1800";
    tmp(59117) := x"1800";
    tmp(59118) := x"2000";
    tmp(59119) := x"2000";
    tmp(59120) := x"2000";
    tmp(59121) := x"2000";
    tmp(59122) := x"2000";
    tmp(59123) := x"2000";
    tmp(59124) := x"2000";
    tmp(59125) := x"2000";
    tmp(59126) := x"1800";
    tmp(59127) := x"1000";
    tmp(59128) := x"0800";
    tmp(59129) := x"1000";
    tmp(59130) := x"1800";
    tmp(59131) := x"2000";
    tmp(59132) := x"2800";
    tmp(59133) := x"2800";
    tmp(59134) := x"2000";
    tmp(59135) := x"2000";
    tmp(59136) := x"2800";
    tmp(59137) := x"2800";
    tmp(59138) := x"3000";
    tmp(59139) := x"2800";
    tmp(59140) := x"3000";
    tmp(59141) := x"3000";
    tmp(59142) := x"3800";
    tmp(59143) := x"4000";
    tmp(59144) := x"4000";
    tmp(59145) := x"4800";
    tmp(59146) := x"4800";
    tmp(59147) := x"4800";
    tmp(59148) := x"4800";
    tmp(59149) := x"5000";
    tmp(59150) := x"5000";
    tmp(59151) := x"5800";
    tmp(59152) := x"5000";
    tmp(59153) := x"5000";
    tmp(59154) := x"4800";
    tmp(59155) := x"3800";
    tmp(59156) := x"3000";
    tmp(59157) := x"3000";
    tmp(59158) := x"4000";
    tmp(59159) := x"4800";
    tmp(59160) := x"4800";
    tmp(59161) := x"4800";
    tmp(59162) := x"4000";
    tmp(59163) := x"4000";
    tmp(59164) := x"5000";
    tmp(59165) := x"6000";
    tmp(59166) := x"6000";
    tmp(59167) := x"6000";
    tmp(59168) := x"5800";
    tmp(59169) := x"5800";
    tmp(59170) := x"6000";
    tmp(59171) := x"6000";
    tmp(59172) := x"6000";
    tmp(59173) := x"6000";
    tmp(59174) := x"6000";
    tmp(59175) := x"6000";
    tmp(59176) := x"6800";
    tmp(59177) := x"5800";
    tmp(59178) := x"6000";
    tmp(59179) := x"7000";
    tmp(59180) := x"6000";
    tmp(59181) := x"5000";
    tmp(59182) := x"5000";
    tmp(59183) := x"5000";
    tmp(59184) := x"5800";
    tmp(59185) := x"5800";
    tmp(59186) := x"6000";
    tmp(59187) := x"5800";
    tmp(59188) := x"6020";
    tmp(59189) := x"7820";
    tmp(59190) := x"7820";
    tmp(59191) := x"6020";
    tmp(59192) := x"7020";
    tmp(59193) := x"7820";
    tmp(59194) := x"8020";
    tmp(59195) := x"7820";
    tmp(59196) := x"7020";
    tmp(59197) := x"8820";
    tmp(59198) := x"8820";
    tmp(59199) := x"8820";
    tmp(59200) := x"8020";
    tmp(59201) := x"9820";
    tmp(59202) := x"9020";
    tmp(59203) := x"8020";
    tmp(59204) := x"5800";
    tmp(59205) := x"6800";
    tmp(59206) := x"7800";
    tmp(59207) := x"9020";
    tmp(59208) := x"b020";
    tmp(59209) := x"e041";
    tmp(59210) := x"f8c3";
    tmp(59211) := x"f9c8";
    tmp(59212) := x"faee";
    tmp(59213) := x"fa4a";
    tmp(59214) := x"f924";
    tmp(59215) := x"f061";
    tmp(59216) := x"f041";
    tmp(59217) := x"a800";
    tmp(59218) := x"d820";
    tmp(59219) := x"f040";
    tmp(59220) := x"d020";
    tmp(59221) := x"d820";
    tmp(59222) := x"a000";
    tmp(59223) := x"9820";
    tmp(59224) := x"3861";
    tmp(59225) := x"0840";
    tmp(59226) := x"0861";
    tmp(59227) := x"1061";
    tmp(59228) := x"0861";
    tmp(59229) := x"1061";
    tmp(59230) := x"1061";
    tmp(59231) := x"1081";
    tmp(59232) := x"1081";
    tmp(59233) := x"10a2";
    tmp(59234) := x"10a2";
    tmp(59235) := x"18c2";
    tmp(59236) := x"18c3";
    tmp(59237) := x"18e3";
    tmp(59238) := x"20e3";
    tmp(59239) := x"2104";
    tmp(59240) := x"2104";
    tmp(59241) := x"2104";
    tmp(59242) := x"2925";
    tmp(59243) := x"2945";
    tmp(59244) := x"2946";
    tmp(59245) := x"2966";
    tmp(59246) := x"2966";
    tmp(59247) := x"3187";
    tmp(59248) := x"3187";
    tmp(59249) := x"3187";
    tmp(59250) := x"31a7";
    tmp(59251) := x"31a8";
    tmp(59252) := x"39c8";
    tmp(59253) := x"39c8";
    tmp(59254) := x"39c8";
    tmp(59255) := x"39c8";
    tmp(59256) := x"39c9";
    tmp(59257) := x"39e9";
    tmp(59258) := x"39c9";
    tmp(59259) := x"39e9";
    tmp(59260) := x"39e9";
    tmp(59261) := x"39e9";
    tmp(59262) := x"39c9";
    tmp(59263) := x"39c8";
    tmp(59264) := x"31a7";
    tmp(59265) := x"2986";
    tmp(59266) := x"2966";
    tmp(59267) := x"2945";
    tmp(59268) := x"2104";
    tmp(59269) := x"18e3";
    tmp(59270) := x"18c3";
    tmp(59271) := x"10c2";
    tmp(59272) := x"10a2";
    tmp(59273) := x"1081";
    tmp(59274) := x"1081";
    tmp(59275) := x"0861";
    tmp(59276) := x"0861";
    tmp(59277) := x"0861";
    tmp(59278) := x"0861";
    tmp(59279) := x"0861";
    tmp(59280) := x"0000";
    tmp(59281) := x"0800";
    tmp(59282) := x"0800";
    tmp(59283) := x"0800";
    tmp(59284) := x"0800";
    tmp(59285) := x"0800";
    tmp(59286) := x"0800";
    tmp(59287) := x"1000";
    tmp(59288) := x"1000";
    tmp(59289) := x"1000";
    tmp(59290) := x"1000";
    tmp(59291) := x"1000";
    tmp(59292) := x"1000";
    tmp(59293) := x"1000";
    tmp(59294) := x"1000";
    tmp(59295) := x"1000";
    tmp(59296) := x"1000";
    tmp(59297) := x"1000";
    tmp(59298) := x"1000";
    tmp(59299) := x"1000";
    tmp(59300) := x"1000";
    tmp(59301) := x"1000";
    tmp(59302) := x"1000";
    tmp(59303) := x"1000";
    tmp(59304) := x"1000";
    tmp(59305) := x"1000";
    tmp(59306) := x"1800";
    tmp(59307) := x"1800";
    tmp(59308) := x"1800";
    tmp(59309) := x"1800";
    tmp(59310) := x"2000";
    tmp(59311) := x"2000";
    tmp(59312) := x"2000";
    tmp(59313) := x"2000";
    tmp(59314) := x"2000";
    tmp(59315) := x"2000";
    tmp(59316) := x"2000";
    tmp(59317) := x"2000";
    tmp(59318) := x"2000";
    tmp(59319) := x"2000";
    tmp(59320) := x"2000";
    tmp(59321) := x"2800";
    tmp(59322) := x"2800";
    tmp(59323) := x"2000";
    tmp(59324) := x"2000";
    tmp(59325) := x"2800";
    tmp(59326) := x"2800";
    tmp(59327) := x"2800";
    tmp(59328) := x"2800";
    tmp(59329) := x"2800";
    tmp(59330) := x"2000";
    tmp(59331) := x"2000";
    tmp(59332) := x"2800";
    tmp(59333) := x"2800";
    tmp(59334) := x"2800";
    tmp(59335) := x"2800";
    tmp(59336) := x"2800";
    tmp(59337) := x"2800";
    tmp(59338) := x"2800";
    tmp(59339) := x"2800";
    tmp(59340) := x"2800";
    tmp(59341) := x"2800";
    tmp(59342) := x"2800";
    tmp(59343) := x"2800";
    tmp(59344) := x"2800";
    tmp(59345) := x"2800";
    tmp(59346) := x"2800";
    tmp(59347) := x"2000";
    tmp(59348) := x"2000";
    tmp(59349) := x"2000";
    tmp(59350) := x"1800";
    tmp(59351) := x"1800";
    tmp(59352) := x"1800";
    tmp(59353) := x"1000";
    tmp(59354) := x"1000";
    tmp(59355) := x"1000";
    tmp(59356) := x"1800";
    tmp(59357) := x"1800";
    tmp(59358) := x"2000";
    tmp(59359) := x"1800";
    tmp(59360) := x"1800";
    tmp(59361) := x"1800";
    tmp(59362) := x"1800";
    tmp(59363) := x"2000";
    tmp(59364) := x"2000";
    tmp(59365) := x"1800";
    tmp(59366) := x"1000";
    tmp(59367) := x"0800";
    tmp(59368) := x"0800";
    tmp(59369) := x"0800";
    tmp(59370) := x"0800";
    tmp(59371) := x"1000";
    tmp(59372) := x"1800";
    tmp(59373) := x"2000";
    tmp(59374) := x"2000";
    tmp(59375) := x"2000";
    tmp(59376) := x"2000";
    tmp(59377) := x"2000";
    tmp(59378) := x"2800";
    tmp(59379) := x"3000";
    tmp(59380) := x"3000";
    tmp(59381) := x"3000";
    tmp(59382) := x"3800";
    tmp(59383) := x"4000";
    tmp(59384) := x"4000";
    tmp(59385) := x"4000";
    tmp(59386) := x"3800";
    tmp(59387) := x"4000";
    tmp(59388) := x"4800";
    tmp(59389) := x"5000";
    tmp(59390) := x"5000";
    tmp(59391) := x"5000";
    tmp(59392) := x"5000";
    tmp(59393) := x"4800";
    tmp(59394) := x"4000";
    tmp(59395) := x"4800";
    tmp(59396) := x"4800";
    tmp(59397) := x"4800";
    tmp(59398) := x"4800";
    tmp(59399) := x"4800";
    tmp(59400) := x"4800";
    tmp(59401) := x"4000";
    tmp(59402) := x"4000";
    tmp(59403) := x"4800";
    tmp(59404) := x"5000";
    tmp(59405) := x"5800";
    tmp(59406) := x"6020";
    tmp(59407) := x"5800";
    tmp(59408) := x"5800";
    tmp(59409) := x"5800";
    tmp(59410) := x"6000";
    tmp(59411) := x"5800";
    tmp(59412) := x"6000";
    tmp(59413) := x"6800";
    tmp(59414) := x"6800";
    tmp(59415) := x"6800";
    tmp(59416) := x"5800";
    tmp(59417) := x"6800";
    tmp(59418) := x"6800";
    tmp(59419) := x"6800";
    tmp(59420) := x"7020";
    tmp(59421) := x"5800";
    tmp(59422) := x"5000";
    tmp(59423) := x"5800";
    tmp(59424) := x"6000";
    tmp(59425) := x"5800";
    tmp(59426) := x"6820";
    tmp(59427) := x"5000";
    tmp(59428) := x"6020";
    tmp(59429) := x"7820";
    tmp(59430) := x"7820";
    tmp(59431) := x"5820";
    tmp(59432) := x"6820";
    tmp(59433) := x"8020";
    tmp(59434) := x"8020";
    tmp(59435) := x"7820";
    tmp(59436) := x"7020";
    tmp(59437) := x"9020";
    tmp(59438) := x"9840";
    tmp(59439) := x"8820";
    tmp(59440) := x"8820";
    tmp(59441) := x"8820";
    tmp(59442) := x"9820";
    tmp(59443) := x"8020";
    tmp(59444) := x"6800";
    tmp(59445) := x"5800";
    tmp(59446) := x"7800";
    tmp(59447) := x"a020";
    tmp(59448) := x"a820";
    tmp(59449) := x"c020";
    tmp(59450) := x"e061";
    tmp(59451) := x"f104";
    tmp(59452) := x"fb2e";
    tmp(59453) := x"fa8b";
    tmp(59454) := x"f924";
    tmp(59455) := x"e881";
    tmp(59456) := x"c820";
    tmp(59457) := x"a800";
    tmp(59458) := x"d020";
    tmp(59459) := x"e020";
    tmp(59460) := x"b820";
    tmp(59461) := x"d020";
    tmp(59462) := x"a020";
    tmp(59463) := x"8041";
    tmp(59464) := x"1841";
    tmp(59465) := x"0861";
    tmp(59466) := x"1061";
    tmp(59467) := x"1061";
    tmp(59468) := x"1061";
    tmp(59469) := x"1081";
    tmp(59470) := x"1081";
    tmp(59471) := x"1082";
    tmp(59472) := x"10a2";
    tmp(59473) := x"10a2";
    tmp(59474) := x"18c2";
    tmp(59475) := x"18c3";
    tmp(59476) := x"20e4";
    tmp(59477) := x"2104";
    tmp(59478) := x"2104";
    tmp(59479) := x"2104";
    tmp(59480) := x"2105";
    tmp(59481) := x"2925";
    tmp(59482) := x"2945";
    tmp(59483) := x"2946";
    tmp(59484) := x"2966";
    tmp(59485) := x"3187";
    tmp(59486) := x"3187";
    tmp(59487) := x"3187";
    tmp(59488) := x"39a8";
    tmp(59489) := x"31a8";
    tmp(59490) := x"39a8";
    tmp(59491) := x"39a8";
    tmp(59492) := x"39a9";
    tmp(59493) := x"39c9";
    tmp(59494) := x"39c9";
    tmp(59495) := x"39c9";
    tmp(59496) := x"39c9";
    tmp(59497) := x"39e9";
    tmp(59498) := x"39ea";
    tmp(59499) := x"39ea";
    tmp(59500) := x"39ea";
    tmp(59501) := x"39ea";
    tmp(59502) := x"39c9";
    tmp(59503) := x"39c9";
    tmp(59504) := x"31a8";
    tmp(59505) := x"3186";
    tmp(59506) := x"2966";
    tmp(59507) := x"2145";
    tmp(59508) := x"2124";
    tmp(59509) := x"18e4";
    tmp(59510) := x"18e3";
    tmp(59511) := x"10c2";
    tmp(59512) := x"10a2";
    tmp(59513) := x"1081";
    tmp(59514) := x"1081";
    tmp(59515) := x"0881";
    tmp(59516) := x"0861";
    tmp(59517) := x"0861";
    tmp(59518) := x"0861";
    tmp(59519) := x"0861";
    tmp(59520) := x"0000";
    tmp(59521) := x"0800";
    tmp(59522) := x"0800";
    tmp(59523) := x"0800";
    tmp(59524) := x"0800";
    tmp(59525) := x"0800";
    tmp(59526) := x"0800";
    tmp(59527) := x"0800";
    tmp(59528) := x"1000";
    tmp(59529) := x"1000";
    tmp(59530) := x"1000";
    tmp(59531) := x"1000";
    tmp(59532) := x"1000";
    tmp(59533) := x"1000";
    tmp(59534) := x"1000";
    tmp(59535) := x"1000";
    tmp(59536) := x"1000";
    tmp(59537) := x"1000";
    tmp(59538) := x"1000";
    tmp(59539) := x"1000";
    tmp(59540) := x"1000";
    tmp(59541) := x"1000";
    tmp(59542) := x"1000";
    tmp(59543) := x"1000";
    tmp(59544) := x"1000";
    tmp(59545) := x"1000";
    tmp(59546) := x"1800";
    tmp(59547) := x"1800";
    tmp(59548) := x"1800";
    tmp(59549) := x"2000";
    tmp(59550) := x"2000";
    tmp(59551) := x"2000";
    tmp(59552) := x"2800";
    tmp(59553) := x"2800";
    tmp(59554) := x"2800";
    tmp(59555) := x"2000";
    tmp(59556) := x"2000";
    tmp(59557) := x"2000";
    tmp(59558) := x"2000";
    tmp(59559) := x"2000";
    tmp(59560) := x"2000";
    tmp(59561) := x"2000";
    tmp(59562) := x"2800";
    tmp(59563) := x"2000";
    tmp(59564) := x"2000";
    tmp(59565) := x"2000";
    tmp(59566) := x"2800";
    tmp(59567) := x"2800";
    tmp(59568) := x"2800";
    tmp(59569) := x"2800";
    tmp(59570) := x"2800";
    tmp(59571) := x"2800";
    tmp(59572) := x"2800";
    tmp(59573) := x"2800";
    tmp(59574) := x"2800";
    tmp(59575) := x"2800";
    tmp(59576) := x"2800";
    tmp(59577) := x"2800";
    tmp(59578) := x"2800";
    tmp(59579) := x"2800";
    tmp(59580) := x"2800";
    tmp(59581) := x"2800";
    tmp(59582) := x"2800";
    tmp(59583) := x"2800";
    tmp(59584) := x"2000";
    tmp(59585) := x"2000";
    tmp(59586) := x"2000";
    tmp(59587) := x"2000";
    tmp(59588) := x"2000";
    tmp(59589) := x"2000";
    tmp(59590) := x"2000";
    tmp(59591) := x"1800";
    tmp(59592) := x"1800";
    tmp(59593) := x"1000";
    tmp(59594) := x"1000";
    tmp(59595) := x"1000";
    tmp(59596) := x"1800";
    tmp(59597) := x"2000";
    tmp(59598) := x"1800";
    tmp(59599) := x"1800";
    tmp(59600) := x"1800";
    tmp(59601) := x"1800";
    tmp(59602) := x"1800";
    tmp(59603) := x"1800";
    tmp(59604) := x"1000";
    tmp(59605) := x"1000";
    tmp(59606) := x"0800";
    tmp(59607) := x"0800";
    tmp(59608) := x"0800";
    tmp(59609) := x"0800";
    tmp(59610) := x"0000";
    tmp(59611) := x"0000";
    tmp(59612) := x"0000";
    tmp(59613) := x"0800";
    tmp(59614) := x"1000";
    tmp(59615) := x"1000";
    tmp(59616) := x"1800";
    tmp(59617) := x"2000";
    tmp(59618) := x"3000";
    tmp(59619) := x"3000";
    tmp(59620) := x"3000";
    tmp(59621) := x"3800";
    tmp(59622) := x"4000";
    tmp(59623) := x"4000";
    tmp(59624) := x"4000";
    tmp(59625) := x"4000";
    tmp(59626) := x"4800";
    tmp(59627) := x"4000";
    tmp(59628) := x"4800";
    tmp(59629) := x"5000";
    tmp(59630) := x"5000";
    tmp(59631) := x"5000";
    tmp(59632) := x"4800";
    tmp(59633) := x"4000";
    tmp(59634) := x"4000";
    tmp(59635) := x"5000";
    tmp(59636) := x"4800";
    tmp(59637) := x"4800";
    tmp(59638) := x"4800";
    tmp(59639) := x"4800";
    tmp(59640) := x"4000";
    tmp(59641) := x"4000";
    tmp(59642) := x"4000";
    tmp(59643) := x"4800";
    tmp(59644) := x"5000";
    tmp(59645) := x"5800";
    tmp(59646) := x"5800";
    tmp(59647) := x"5000";
    tmp(59648) := x"5800";
    tmp(59649) := x"5800";
    tmp(59650) := x"5800";
    tmp(59651) := x"5800";
    tmp(59652) := x"6000";
    tmp(59653) := x"6000";
    tmp(59654) := x"6800";
    tmp(59655) := x"6800";
    tmp(59656) := x"6000";
    tmp(59657) := x"8820";
    tmp(59658) := x"7820";
    tmp(59659) := x"7020";
    tmp(59660) := x"7820";
    tmp(59661) := x"6020";
    tmp(59662) := x"5800";
    tmp(59663) := x"5800";
    tmp(59664) := x"6000";
    tmp(59665) := x"5800";
    tmp(59666) := x"6820";
    tmp(59667) := x"6000";
    tmp(59668) := x"7020";
    tmp(59669) := x"7820";
    tmp(59670) := x"7820";
    tmp(59671) := x"6820";
    tmp(59672) := x"6820";
    tmp(59673) := x"8020";
    tmp(59674) := x"8820";
    tmp(59675) := x"8020";
    tmp(59676) := x"7820";
    tmp(59677) := x"8820";
    tmp(59678) := x"a840";
    tmp(59679) := x"8020";
    tmp(59680) := x"8820";
    tmp(59681) := x"8020";
    tmp(59682) := x"9020";
    tmp(59683) := x"8020";
    tmp(59684) := x"7820";
    tmp(59685) := x"5800";
    tmp(59686) := x"7000";
    tmp(59687) := x"9820";
    tmp(59688) := x"b020";
    tmp(59689) := x"a820";
    tmp(59690) := x"c820";
    tmp(59691) := x"e041";
    tmp(59692) := x"f0e3";
    tmp(59693) := x"e925";
    tmp(59694) := x"f0e3";
    tmp(59695) := x"e861";
    tmp(59696) := x"c820";
    tmp(59697) := x"a800";
    tmp(59698) := x"c820";
    tmp(59699) := x"d020";
    tmp(59700) := x"b020";
    tmp(59701) := x"c820";
    tmp(59702) := x"a020";
    tmp(59703) := x"5841";
    tmp(59704) := x"1041";
    tmp(59705) := x"1061";
    tmp(59706) := x"1061";
    tmp(59707) := x"1061";
    tmp(59708) := x"1081";
    tmp(59709) := x"1081";
    tmp(59710) := x"10a2";
    tmp(59711) := x"18a2";
    tmp(59712) := x"18c2";
    tmp(59713) := x"18c3";
    tmp(59714) := x"18e3";
    tmp(59715) := x"20e3";
    tmp(59716) := x"18e3";
    tmp(59717) := x"2104";
    tmp(59718) := x"2104";
    tmp(59719) := x"2925";
    tmp(59720) := x"2925";
    tmp(59721) := x"2945";
    tmp(59722) := x"2966";
    tmp(59723) := x"3186";
    tmp(59724) := x"3187";
    tmp(59725) := x"3187";
    tmp(59726) := x"3187";
    tmp(59727) := x"39a8";
    tmp(59728) := x"39a8";
    tmp(59729) := x"39c8";
    tmp(59730) := x"39c8";
    tmp(59731) := x"39e9";
    tmp(59732) := x"39c8";
    tmp(59733) := x"39c9";
    tmp(59734) := x"39c9";
    tmp(59735) := x"39c9";
    tmp(59736) := x"39c9";
    tmp(59737) := x"39e9";
    tmp(59738) := x"39c9";
    tmp(59739) := x"39c9";
    tmp(59740) := x"39a9";
    tmp(59741) := x"31a9";
    tmp(59742) := x"31a9";
    tmp(59743) := x"31a9";
    tmp(59744) := x"3188";
    tmp(59745) := x"3187";
    tmp(59746) := x"2966";
    tmp(59747) := x"2145";
    tmp(59748) := x"2104";
    tmp(59749) := x"18e4";
    tmp(59750) := x"18c3";
    tmp(59751) := x"10c2";
    tmp(59752) := x"10a2";
    tmp(59753) := x"1081";
    tmp(59754) := x"1081";
    tmp(59755) := x"0861";
    tmp(59756) := x"0861";
    tmp(59757) := x"0861";
    tmp(59758) := x"0861";
    tmp(59759) := x"0861";
    tmp(59760) := x"0000";
    tmp(59761) := x"0800";
    tmp(59762) := x"0800";
    tmp(59763) := x"0800";
    tmp(59764) := x"0800";
    tmp(59765) := x"0800";
    tmp(59766) := x"0800";
    tmp(59767) := x"0800";
    tmp(59768) := x"0800";
    tmp(59769) := x"1000";
    tmp(59770) := x"1000";
    tmp(59771) := x"1000";
    tmp(59772) := x"1000";
    tmp(59773) := x"1000";
    tmp(59774) := x"1000";
    tmp(59775) := x"1000";
    tmp(59776) := x"1000";
    tmp(59777) := x"1000";
    tmp(59778) := x"1000";
    tmp(59779) := x"1000";
    tmp(59780) := x"1000";
    tmp(59781) := x"1000";
    tmp(59782) := x"1000";
    tmp(59783) := x"1000";
    tmp(59784) := x"1000";
    tmp(59785) := x"1000";
    tmp(59786) := x"1800";
    tmp(59787) := x"1800";
    tmp(59788) := x"2000";
    tmp(59789) := x"2000";
    tmp(59790) := x"2000";
    tmp(59791) := x"2000";
    tmp(59792) := x"2800";
    tmp(59793) := x"2800";
    tmp(59794) := x"2000";
    tmp(59795) := x"2000";
    tmp(59796) := x"2000";
    tmp(59797) := x"2800";
    tmp(59798) := x"2800";
    tmp(59799) := x"2000";
    tmp(59800) := x"2000";
    tmp(59801) := x"2000";
    tmp(59802) := x"2000";
    tmp(59803) := x"2000";
    tmp(59804) := x"2000";
    tmp(59805) := x"2000";
    tmp(59806) := x"2800";
    tmp(59807) := x"2800";
    tmp(59808) := x"2800";
    tmp(59809) := x"2800";
    tmp(59810) := x"2800";
    tmp(59811) := x"2800";
    tmp(59812) := x"2800";
    tmp(59813) := x"2800";
    tmp(59814) := x"2800";
    tmp(59815) := x"2800";
    tmp(59816) := x"2800";
    tmp(59817) := x"2800";
    tmp(59818) := x"2800";
    tmp(59819) := x"2800";
    tmp(59820) := x"2800";
    tmp(59821) := x"2800";
    tmp(59822) := x"2800";
    tmp(59823) := x"2000";
    tmp(59824) := x"2000";
    tmp(59825) := x"2000";
    tmp(59826) := x"2000";
    tmp(59827) := x"2000";
    tmp(59828) := x"2000";
    tmp(59829) := x"2000";
    tmp(59830) := x"2000";
    tmp(59831) := x"1800";
    tmp(59832) := x"1800";
    tmp(59833) := x"1000";
    tmp(59834) := x"1000";
    tmp(59835) := x"1800";
    tmp(59836) := x"1800";
    tmp(59837) := x"1800";
    tmp(59838) := x"1800";
    tmp(59839) := x"1800";
    tmp(59840) := x"1800";
    tmp(59841) := x"1800";
    tmp(59842) := x"1800";
    tmp(59843) := x"1800";
    tmp(59844) := x"1800";
    tmp(59845) := x"1000";
    tmp(59846) := x"1000";
    tmp(59847) := x"1000";
    tmp(59848) := x"0800";
    tmp(59849) := x"0800";
    tmp(59850) := x"0800";
    tmp(59851) := x"1000";
    tmp(59852) := x"1000";
    tmp(59853) := x"1000";
    tmp(59854) := x"1000";
    tmp(59855) := x"1000";
    tmp(59856) := x"1800";
    tmp(59857) := x"2800";
    tmp(59858) := x"3000";
    tmp(59859) := x"3000";
    tmp(59860) := x"3800";
    tmp(59861) := x"4000";
    tmp(59862) := x"4800";
    tmp(59863) := x"4800";
    tmp(59864) := x"4000";
    tmp(59865) := x"4000";
    tmp(59866) := x"4000";
    tmp(59867) := x"4000";
    tmp(59868) := x"5000";
    tmp(59869) := x"5000";
    tmp(59870) := x"5800";
    tmp(59871) := x"5000";
    tmp(59872) := x"4000";
    tmp(59873) := x"4000";
    tmp(59874) := x"4800";
    tmp(59875) := x"5000";
    tmp(59876) := x"5000";
    tmp(59877) := x"4800";
    tmp(59878) := x"5000";
    tmp(59879) := x"4800";
    tmp(59880) := x"4000";
    tmp(59881) := x"4000";
    tmp(59882) := x"4800";
    tmp(59883) := x"4000";
    tmp(59884) := x"4800";
    tmp(59885) := x"5000";
    tmp(59886) := x"5000";
    tmp(59887) := x"5800";
    tmp(59888) := x"5800";
    tmp(59889) := x"5800";
    tmp(59890) := x"5800";
    tmp(59891) := x"5800";
    tmp(59892) := x"5800";
    tmp(59893) := x"6800";
    tmp(59894) := x"7000";
    tmp(59895) := x"6800";
    tmp(59896) := x"7800";
    tmp(59897) := x"8820";
    tmp(59898) := x"7820";
    tmp(59899) := x"8020";
    tmp(59900) := x"7820";
    tmp(59901) := x"6820";
    tmp(59902) := x"5800";
    tmp(59903) := x"5800";
    tmp(59904) := x"6000";
    tmp(59905) := x"5800";
    tmp(59906) := x"6000";
    tmp(59907) := x"6000";
    tmp(59908) := x"6820";
    tmp(59909) := x"8020";
    tmp(59910) := x"6820";
    tmp(59911) := x"7820";
    tmp(59912) := x"6820";
    tmp(59913) := x"7020";
    tmp(59914) := x"8820";
    tmp(59915) := x"8020";
    tmp(59916) := x"7020";
    tmp(59917) := x"8820";
    tmp(59918) := x"9820";
    tmp(59919) := x"8820";
    tmp(59920) := x"8020";
    tmp(59921) := x"8820";
    tmp(59922) := x"9020";
    tmp(59923) := x"8820";
    tmp(59924) := x"8820";
    tmp(59925) := x"6800";
    tmp(59926) := x"7000";
    tmp(59927) := x"8820";
    tmp(59928) := x"b020";
    tmp(59929) := x"a820";
    tmp(59930) := x"c820";
    tmp(59931) := x"d020";
    tmp(59932) := x"e841";
    tmp(59933) := x"d861";
    tmp(59934) := x"e8a2";
    tmp(59935) := x"e861";
    tmp(59936) := x"c820";
    tmp(59937) := x"a800";
    tmp(59938) := x"d820";
    tmp(59939) := x"d820";
    tmp(59940) := x"a800";
    tmp(59941) := x"a820";
    tmp(59942) := x"9820";
    tmp(59943) := x"3861";
    tmp(59944) := x"1061";
    tmp(59945) := x"1061";
    tmp(59946) := x"1081";
    tmp(59947) := x"1081";
    tmp(59948) := x"10a2";
    tmp(59949) := x"10a2";
    tmp(59950) := x"18c2";
    tmp(59951) := x"18c3";
    tmp(59952) := x"18e3";
    tmp(59953) := x"20e4";
    tmp(59954) := x"2104";
    tmp(59955) := x"2104";
    tmp(59956) := x"2124";
    tmp(59957) := x"2104";
    tmp(59958) := x"2125";
    tmp(59959) := x"2925";
    tmp(59960) := x"2945";
    tmp(59961) := x"2966";
    tmp(59962) := x"3186";
    tmp(59963) := x"3187";
    tmp(59964) := x"3187";
    tmp(59965) := x"3187";
    tmp(59966) := x"39a8";
    tmp(59967) := x"31a8";
    tmp(59968) := x"39c8";
    tmp(59969) := x"39a8";
    tmp(59970) := x"39a8";
    tmp(59971) := x"31a8";
    tmp(59972) := x"39a8";
    tmp(59973) := x"39a8";
    tmp(59974) := x"39c9";
    tmp(59975) := x"39a9";
    tmp(59976) := x"31a8";
    tmp(59977) := x"31a8";
    tmp(59978) := x"39a8";
    tmp(59979) := x"39a8";
    tmp(59980) := x"3188";
    tmp(59981) := x"31a8";
    tmp(59982) := x"3188";
    tmp(59983) := x"3188";
    tmp(59984) := x"3188";
    tmp(59985) := x"2967";
    tmp(59986) := x"2946";
    tmp(59987) := x"2145";
    tmp(59988) := x"2124";
    tmp(59989) := x"18e4";
    tmp(59990) := x"18e3";
    tmp(59991) := x"10c3";
    tmp(59992) := x"10a2";
    tmp(59993) := x"10a2";
    tmp(59994) := x"1081";
    tmp(59995) := x"1081";
    tmp(59996) := x"1081";
    tmp(59997) := x"0881";
    tmp(59998) := x"0881";
    tmp(59999) := x"0881";
    tmp(60000) := x"0000";
    tmp(60001) := x"0800";
    tmp(60002) := x"0800";
    tmp(60003) := x"0800";
    tmp(60004) := x"0800";
    tmp(60005) := x"0800";
    tmp(60006) := x"0800";
    tmp(60007) := x"0800";
    tmp(60008) := x"0800";
    tmp(60009) := x"1000";
    tmp(60010) := x"1000";
    tmp(60011) := x"1000";
    tmp(60012) := x"1000";
    tmp(60013) := x"1000";
    tmp(60014) := x"1000";
    tmp(60015) := x"1000";
    tmp(60016) := x"1000";
    tmp(60017) := x"1000";
    tmp(60018) := x"1000";
    tmp(60019) := x"1000";
    tmp(60020) := x"1000";
    tmp(60021) := x"1000";
    tmp(60022) := x"1000";
    tmp(60023) := x"1000";
    tmp(60024) := x"1000";
    tmp(60025) := x"1800";
    tmp(60026) := x"1800";
    tmp(60027) := x"2000";
    tmp(60028) := x"2000";
    tmp(60029) := x"2000";
    tmp(60030) := x"2000";
    tmp(60031) := x"2800";
    tmp(60032) := x"2800";
    tmp(60033) := x"2000";
    tmp(60034) := x"2000";
    tmp(60035) := x"2000";
    tmp(60036) := x"2800";
    tmp(60037) := x"2000";
    tmp(60038) := x"2000";
    tmp(60039) := x"2800";
    tmp(60040) := x"2000";
    tmp(60041) := x"2000";
    tmp(60042) := x"2000";
    tmp(60043) := x"2000";
    tmp(60044) := x"2000";
    tmp(60045) := x"2800";
    tmp(60046) := x"2800";
    tmp(60047) := x"2800";
    tmp(60048) := x"2800";
    tmp(60049) := x"2800";
    tmp(60050) := x"2000";
    tmp(60051) := x"2000";
    tmp(60052) := x"2000";
    tmp(60053) := x"2000";
    tmp(60054) := x"2000";
    tmp(60055) := x"2800";
    tmp(60056) := x"2800";
    tmp(60057) := x"2800";
    tmp(60058) := x"2800";
    tmp(60059) := x"2800";
    tmp(60060) := x"2800";
    tmp(60061) := x"2000";
    tmp(60062) := x"2000";
    tmp(60063) := x"2000";
    tmp(60064) := x"2000";
    tmp(60065) := x"2000";
    tmp(60066) := x"2000";
    tmp(60067) := x"2000";
    tmp(60068) := x"2000";
    tmp(60069) := x"2000";
    tmp(60070) := x"2000";
    tmp(60071) := x"1800";
    tmp(60072) := x"1800";
    tmp(60073) := x"1800";
    tmp(60074) := x"2000";
    tmp(60075) := x"1800";
    tmp(60076) := x"1000";
    tmp(60077) := x"1800";
    tmp(60078) := x"2000";
    tmp(60079) := x"2000";
    tmp(60080) := x"2000";
    tmp(60081) := x"2000";
    tmp(60082) := x"2000";
    tmp(60083) := x"2000";
    tmp(60084) := x"2000";
    tmp(60085) := x"1800";
    tmp(60086) := x"1000";
    tmp(60087) := x"1000";
    tmp(60088) := x"1000";
    tmp(60089) := x"1800";
    tmp(60090) := x"1800";
    tmp(60091) := x"1800";
    tmp(60092) := x"1800";
    tmp(60093) := x"1800";
    tmp(60094) := x"1800";
    tmp(60095) := x"1800";
    tmp(60096) := x"2000";
    tmp(60097) := x"2800";
    tmp(60098) := x"3000";
    tmp(60099) := x"3000";
    tmp(60100) := x"3800";
    tmp(60101) := x"4000";
    tmp(60102) := x"4000";
    tmp(60103) := x"4000";
    tmp(60104) := x"4000";
    tmp(60105) := x"4000";
    tmp(60106) := x"4000";
    tmp(60107) := x"4800";
    tmp(60108) := x"4800";
    tmp(60109) := x"5000";
    tmp(60110) := x"5000";
    tmp(60111) := x"5000";
    tmp(60112) := x"5000";
    tmp(60113) := x"5000";
    tmp(60114) := x"5000";
    tmp(60115) := x"5000";
    tmp(60116) := x"5000";
    tmp(60117) := x"5000";
    tmp(60118) := x"5000";
    tmp(60119) := x"4800";
    tmp(60120) := x"4000";
    tmp(60121) := x"4000";
    tmp(60122) := x"4000";
    tmp(60123) := x"4000";
    tmp(60124) := x"5000";
    tmp(60125) := x"5800";
    tmp(60126) := x"5800";
    tmp(60127) := x"5800";
    tmp(60128) := x"5800";
    tmp(60129) := x"5000";
    tmp(60130) := x"5000";
    tmp(60131) := x"5000";
    tmp(60132) := x"6000";
    tmp(60133) := x"7000";
    tmp(60134) := x"6800";
    tmp(60135) := x"6800";
    tmp(60136) := x"7800";
    tmp(60137) := x"7000";
    tmp(60138) := x"7820";
    tmp(60139) := x"8020";
    tmp(60140) := x"8020";
    tmp(60141) := x"6820";
    tmp(60142) := x"6820";
    tmp(60143) := x"6020";
    tmp(60144) := x"5800";
    tmp(60145) := x"5800";
    tmp(60146) := x"5800";
    tmp(60147) := x"6000";
    tmp(60148) := x"6000";
    tmp(60149) := x"9040";
    tmp(60150) := x"6820";
    tmp(60151) := x"7020";
    tmp(60152) := x"7020";
    tmp(60153) := x"7020";
    tmp(60154) := x"8020";
    tmp(60155) := x"9040";
    tmp(60156) := x"7020";
    tmp(60157) := x"8820";
    tmp(60158) := x"a020";
    tmp(60159) := x"8820";
    tmp(60160) := x"7820";
    tmp(60161) := x"9020";
    tmp(60162) := x"9020";
    tmp(60163) := x"8820";
    tmp(60164) := x"9820";
    tmp(60165) := x"6800";
    tmp(60166) := x"6800";
    tmp(60167) := x"8000";
    tmp(60168) := x"a020";
    tmp(60169) := x"b020";
    tmp(60170) := x"c820";
    tmp(60171) := x"d820";
    tmp(60172) := x"d820";
    tmp(60173) := x"c020";
    tmp(60174) := x"e061";
    tmp(60175) := x"e841";
    tmp(60176) := x"c820";
    tmp(60177) := x"b000";
    tmp(60178) := x"c020";
    tmp(60179) := x"c020";
    tmp(60180) := x"9800";
    tmp(60181) := x"9820";
    tmp(60182) := x"8020";
    tmp(60183) := x"2061";
    tmp(60184) := x"1061";
    tmp(60185) := x"1081";
    tmp(60186) := x"1081";
    tmp(60187) := x"10a2";
    tmp(60188) := x"18a2";
    tmp(60189) := x"18c2";
    tmp(60190) := x"18c3";
    tmp(60191) := x"18e3";
    tmp(60192) := x"20e4";
    tmp(60193) := x"2104";
    tmp(60194) := x"2104";
    tmp(60195) := x"2125";
    tmp(60196) := x"2125";
    tmp(60197) := x"2925";
    tmp(60198) := x"2945";
    tmp(60199) := x"2946";
    tmp(60200) := x"2966";
    tmp(60201) := x"3166";
    tmp(60202) := x"3187";
    tmp(60203) := x"3187";
    tmp(60204) := x"3187";
    tmp(60205) := x"31a7";
    tmp(60206) := x"31a8";
    tmp(60207) := x"39a8";
    tmp(60208) := x"31a8";
    tmp(60209) := x"39a8";
    tmp(60210) := x"31a8";
    tmp(60211) := x"31a8";
    tmp(60212) := x"31a8";
    tmp(60213) := x"3188";
    tmp(60214) := x"3188";
    tmp(60215) := x"31a8";
    tmp(60216) := x"31a9";
    tmp(60217) := x"31a8";
    tmp(60218) := x"31a8";
    tmp(60219) := x"31a8";
    tmp(60220) := x"3187";
    tmp(60221) := x"3187";
    tmp(60222) := x"2987";
    tmp(60223) := x"3187";
    tmp(60224) := x"2987";
    tmp(60225) := x"2967";
    tmp(60226) := x"2946";
    tmp(60227) := x"2125";
    tmp(60228) := x"2104";
    tmp(60229) := x"1904";
    tmp(60230) := x"1903";
    tmp(60231) := x"18e3";
    tmp(60232) := x"18c3";
    tmp(60233) := x"10c2";
    tmp(60234) := x"10c2";
    tmp(60235) := x"10c2";
    tmp(60236) := x"10a2";
    tmp(60237) := x"10a2";
    tmp(60238) := x"10a2";
    tmp(60239) := x"10a2";
    tmp(60240) := x"0000";
    tmp(60241) := x"0800";
    tmp(60242) := x"0800";
    tmp(60243) := x"0800";
    tmp(60244) := x"0800";
    tmp(60245) := x"0800";
    tmp(60246) := x"0800";
    tmp(60247) := x"0800";
    tmp(60248) := x"0800";
    tmp(60249) := x"0800";
    tmp(60250) := x"0800";
    tmp(60251) := x"1000";
    tmp(60252) := x"1000";
    tmp(60253) := x"1000";
    tmp(60254) := x"1000";
    tmp(60255) := x"1000";
    tmp(60256) := x"1000";
    tmp(60257) := x"1000";
    tmp(60258) := x"1000";
    tmp(60259) := x"1000";
    tmp(60260) := x"1000";
    tmp(60261) := x"1000";
    tmp(60262) := x"1000";
    tmp(60263) := x"1000";
    tmp(60264) := x"1800";
    tmp(60265) := x"1800";
    tmp(60266) := x"1800";
    tmp(60267) := x"2000";
    tmp(60268) := x"2000";
    tmp(60269) := x"2000";
    tmp(60270) := x"2000";
    tmp(60271) := x"2000";
    tmp(60272) := x"2000";
    tmp(60273) := x"2000";
    tmp(60274) := x"2000";
    tmp(60275) := x"2000";
    tmp(60276) := x"2000";
    tmp(60277) := x"1800";
    tmp(60278) := x"1800";
    tmp(60279) := x"2000";
    tmp(60280) := x"2000";
    tmp(60281) := x"2000";
    tmp(60282) := x"2000";
    tmp(60283) := x"2000";
    tmp(60284) := x"2000";
    tmp(60285) := x"2000";
    tmp(60286) := x"2800";
    tmp(60287) := x"2800";
    tmp(60288) := x"2800";
    tmp(60289) := x"2800";
    tmp(60290) := x"2800";
    tmp(60291) := x"2800";
    tmp(60292) := x"2800";
    tmp(60293) := x"2000";
    tmp(60294) := x"2000";
    tmp(60295) := x"2800";
    tmp(60296) := x"2800";
    tmp(60297) := x"2800";
    tmp(60298) := x"2800";
    tmp(60299) := x"2000";
    tmp(60300) := x"2000";
    tmp(60301) := x"2000";
    tmp(60302) := x"2000";
    tmp(60303) := x"2000";
    tmp(60304) := x"2800";
    tmp(60305) := x"2800";
    tmp(60306) := x"2800";
    tmp(60307) := x"2800";
    tmp(60308) := x"2000";
    tmp(60309) := x"2000";
    tmp(60310) := x"2000";
    tmp(60311) := x"2000";
    tmp(60312) := x"2000";
    tmp(60313) := x"2000";
    tmp(60314) := x"1000";
    tmp(60315) := x"1000";
    tmp(60316) := x"1800";
    tmp(60317) := x"2000";
    tmp(60318) := x"2000";
    tmp(60319) := x"2000";
    tmp(60320) := x"2000";
    tmp(60321) := x"2000";
    tmp(60322) := x"2000";
    tmp(60323) := x"2000";
    tmp(60324) := x"2000";
    tmp(60325) := x"1800";
    tmp(60326) := x"1000";
    tmp(60327) := x"1000";
    tmp(60328) := x"1000";
    tmp(60329) := x"1000";
    tmp(60330) := x"1000";
    tmp(60331) := x"1000";
    tmp(60332) := x"1000";
    tmp(60333) := x"1000";
    tmp(60334) := x"1800";
    tmp(60335) := x"1800";
    tmp(60336) := x"2000";
    tmp(60337) := x"2000";
    tmp(60338) := x"3000";
    tmp(60339) := x"3000";
    tmp(60340) := x"3000";
    tmp(60341) := x"3800";
    tmp(60342) := x"3800";
    tmp(60343) := x"4000";
    tmp(60344) := x"4000";
    tmp(60345) := x"3800";
    tmp(60346) := x"3800";
    tmp(60347) := x"4000";
    tmp(60348) := x"4800";
    tmp(60349) := x"5000";
    tmp(60350) := x"5000";
    tmp(60351) := x"5000";
    tmp(60352) := x"5000";
    tmp(60353) := x"5000";
    tmp(60354) := x"5000";
    tmp(60355) := x"5800";
    tmp(60356) := x"5000";
    tmp(60357) := x"5000";
    tmp(60358) := x"4800";
    tmp(60359) := x"4000";
    tmp(60360) := x"4800";
    tmp(60361) := x"4800";
    tmp(60362) := x"5000";
    tmp(60363) := x"5000";
    tmp(60364) := x"5800";
    tmp(60365) := x"5800";
    tmp(60366) := x"6000";
    tmp(60367) := x"6800";
    tmp(60368) := x"5000";
    tmp(60369) := x"5000";
    tmp(60370) := x"5000";
    tmp(60371) := x"5800";
    tmp(60372) := x"6000";
    tmp(60373) := x"7000";
    tmp(60374) := x"6000";
    tmp(60375) := x"6800";
    tmp(60376) := x"7800";
    tmp(60377) := x"7000";
    tmp(60378) := x"7800";
    tmp(60379) := x"7820";
    tmp(60380) := x"7820";
    tmp(60381) := x"6820";
    tmp(60382) := x"7020";
    tmp(60383) := x"6820";
    tmp(60384) := x"5800";
    tmp(60385) := x"5800";
    tmp(60386) := x"5800";
    tmp(60387) := x"6820";
    tmp(60388) := x"5800";
    tmp(60389) := x"9040";
    tmp(60390) := x"6820";
    tmp(60391) := x"7020";
    tmp(60392) := x"7020";
    tmp(60393) := x"6820";
    tmp(60394) := x"7820";
    tmp(60395) := x"9040";
    tmp(60396) := x"7820";
    tmp(60397) := x"8820";
    tmp(60398) := x"9020";
    tmp(60399) := x"8020";
    tmp(60400) := x"8020";
    tmp(60401) := x"9020";
    tmp(60402) := x"9020";
    tmp(60403) := x"8020";
    tmp(60404) := x"9820";
    tmp(60405) := x"7000";
    tmp(60406) := x"6000";
    tmp(60407) := x"8000";
    tmp(60408) := x"a020";
    tmp(60409) := x"b820";
    tmp(60410) := x"c020";
    tmp(60411) := x"b820";
    tmp(60412) := x"c820";
    tmp(60413) := x"c020";
    tmp(60414) := x"d841";
    tmp(60415) := x"c820";
    tmp(60416) := x"b000";
    tmp(60417) := x"b800";
    tmp(60418) := x"c820";
    tmp(60419) := x"b820";
    tmp(60420) := x"9800";
    tmp(60421) := x"a820";
    tmp(60422) := x"6841";
    tmp(60423) := x"1861";
    tmp(60424) := x"1081";
    tmp(60425) := x"1081";
    tmp(60426) := x"10a2";
    tmp(60427) := x"10a2";
    tmp(60428) := x"18c2";
    tmp(60429) := x"18c3";
    tmp(60430) := x"20e3";
    tmp(60431) := x"20e4";
    tmp(60432) := x"2104";
    tmp(60433) := x"2105";
    tmp(60434) := x"2925";
    tmp(60435) := x"2925";
    tmp(60436) := x"2925";
    tmp(60437) := x"2946";
    tmp(60438) := x"2945";
    tmp(60439) := x"2966";
    tmp(60440) := x"3166";
    tmp(60441) := x"3166";
    tmp(60442) := x"3187";
    tmp(60443) := x"3187";
    tmp(60444) := x"3187";
    tmp(60445) := x"3187";
    tmp(60446) := x"31a8";
    tmp(60447) := x"3187";
    tmp(60448) := x"3187";
    tmp(60449) := x"3188";
    tmp(60450) := x"31a8";
    tmp(60451) := x"3187";
    tmp(60452) := x"3187";
    tmp(60453) := x"3188";
    tmp(60454) := x"3188";
    tmp(60455) := x"3188";
    tmp(60456) := x"3188";
    tmp(60457) := x"3188";
    tmp(60458) := x"3188";
    tmp(60459) := x"3187";
    tmp(60460) := x"2967";
    tmp(60461) := x"2967";
    tmp(60462) := x"2967";
    tmp(60463) := x"2967";
    tmp(60464) := x"2967";
    tmp(60465) := x"2986";
    tmp(60466) := x"2966";
    tmp(60467) := x"2946";
    tmp(60468) := x"2946";
    tmp(60469) := x"2145";
    tmp(60470) := x"2125";
    tmp(60471) := x"2124";
    tmp(60472) := x"2104";
    tmp(60473) := x"1903";
    tmp(60474) := x"1903";
    tmp(60475) := x"18e3";
    tmp(60476) := x"18e3";
    tmp(60477) := x"18e2";
    tmp(60478) := x"18e2";
    tmp(60479) := x"10c2";
    tmp(60480) := x"0000";
    tmp(60481) := x"0800";
    tmp(60482) := x"0800";
    tmp(60483) := x"0800";
    tmp(60484) := x"0800";
    tmp(60485) := x"0800";
    tmp(60486) := x"0800";
    tmp(60487) := x"0800";
    tmp(60488) := x"0800";
    tmp(60489) := x"0800";
    tmp(60490) := x"0800";
    tmp(60491) := x"1000";
    tmp(60492) := x"1000";
    tmp(60493) := x"1000";
    tmp(60494) := x"1000";
    tmp(60495) := x"1000";
    tmp(60496) := x"1000";
    tmp(60497) := x"1000";
    tmp(60498) := x"1000";
    tmp(60499) := x"1000";
    tmp(60500) := x"1000";
    tmp(60501) := x"1800";
    tmp(60502) := x"1800";
    tmp(60503) := x"1800";
    tmp(60504) := x"1000";
    tmp(60505) := x"1800";
    tmp(60506) := x"1800";
    tmp(60507) := x"1800";
    tmp(60508) := x"1800";
    tmp(60509) := x"1800";
    tmp(60510) := x"1800";
    tmp(60511) := x"2000";
    tmp(60512) := x"2000";
    tmp(60513) := x"2000";
    tmp(60514) := x"2000";
    tmp(60515) := x"2000";
    tmp(60516) := x"1800";
    tmp(60517) := x"2000";
    tmp(60518) := x"2000";
    tmp(60519) := x"2000";
    tmp(60520) := x"2000";
    tmp(60521) := x"2000";
    tmp(60522) := x"2000";
    tmp(60523) := x"2000";
    tmp(60524) := x"2000";
    tmp(60525) := x"2000";
    tmp(60526) := x"2000";
    tmp(60527) := x"2000";
    tmp(60528) := x"2000";
    tmp(60529) := x"2000";
    tmp(60530) := x"2800";
    tmp(60531) := x"2800";
    tmp(60532) := x"2800";
    tmp(60533) := x"2800";
    tmp(60534) := x"2800";
    tmp(60535) := x"2000";
    tmp(60536) := x"2000";
    tmp(60537) := x"2000";
    tmp(60538) := x"2000";
    tmp(60539) := x"2800";
    tmp(60540) := x"2800";
    tmp(60541) := x"2000";
    tmp(60542) := x"2000";
    tmp(60543) := x"2800";
    tmp(60544) := x"2800";
    tmp(60545) := x"2800";
    tmp(60546) := x"2800";
    tmp(60547) := x"2800";
    tmp(60548) := x"2800";
    tmp(60549) := x"2000";
    tmp(60550) := x"2000";
    tmp(60551) := x"2000";
    tmp(60552) := x"1800";
    tmp(60553) := x"1000";
    tmp(60554) := x"1000";
    tmp(60555) := x"1000";
    tmp(60556) := x"2000";
    tmp(60557) := x"2000";
    tmp(60558) := x"2000";
    tmp(60559) := x"2000";
    tmp(60560) := x"2000";
    tmp(60561) := x"2000";
    tmp(60562) := x"2800";
    tmp(60563) := x"2000";
    tmp(60564) := x"2000";
    tmp(60565) := x"1800";
    tmp(60566) := x"1000";
    tmp(60567) := x"1000";
    tmp(60568) := x"1000";
    tmp(60569) := x"1000";
    tmp(60570) := x"1000";
    tmp(60571) := x"1000";
    tmp(60572) := x"1000";
    tmp(60573) := x"1000";
    tmp(60574) := x"1000";
    tmp(60575) := x"1000";
    tmp(60576) := x"1800";
    tmp(60577) := x"2000";
    tmp(60578) := x"2800";
    tmp(60579) := x"2800";
    tmp(60580) := x"3000";
    tmp(60581) := x"3800";
    tmp(60582) := x"3800";
    tmp(60583) := x"4000";
    tmp(60584) := x"4000";
    tmp(60585) := x"3800";
    tmp(60586) := x"4000";
    tmp(60587) := x"4000";
    tmp(60588) := x"4800";
    tmp(60589) := x"5000";
    tmp(60590) := x"5000";
    tmp(60591) := x"5000";
    tmp(60592) := x"5000";
    tmp(60593) := x"5000";
    tmp(60594) := x"5000";
    tmp(60595) := x"5800";
    tmp(60596) := x"5000";
    tmp(60597) := x"5000";
    tmp(60598) := x"4800";
    tmp(60599) := x"4000";
    tmp(60600) := x"4800";
    tmp(60601) := x"4800";
    tmp(60602) := x"5000";
    tmp(60603) := x"4800";
    tmp(60604) := x"5000";
    tmp(60605) := x"5800";
    tmp(60606) := x"6000";
    tmp(60607) := x"5800";
    tmp(60608) := x"5000";
    tmp(60609) := x"5000";
    tmp(60610) := x"5000";
    tmp(60611) := x"5800";
    tmp(60612) := x"6800";
    tmp(60613) := x"6800";
    tmp(60614) := x"5800";
    tmp(60615) := x"6000";
    tmp(60616) := x"7000";
    tmp(60617) := x"7000";
    tmp(60618) := x"7800";
    tmp(60619) := x"7820";
    tmp(60620) := x"8820";
    tmp(60621) := x"6800";
    tmp(60622) := x"6820";
    tmp(60623) := x"6820";
    tmp(60624) := x"6020";
    tmp(60625) := x"6820";
    tmp(60626) := x"5800";
    tmp(60627) := x"6820";
    tmp(60628) := x"6000";
    tmp(60629) := x"8820";
    tmp(60630) := x"7820";
    tmp(60631) := x"6820";
    tmp(60632) := x"6820";
    tmp(60633) := x"6020";
    tmp(60634) := x"7020";
    tmp(60635) := x"9020";
    tmp(60636) := x"8820";
    tmp(60637) := x"8020";
    tmp(60638) := x"9020";
    tmp(60639) := x"8020";
    tmp(60640) := x"8820";
    tmp(60641) := x"8820";
    tmp(60642) := x"9820";
    tmp(60643) := x"8820";
    tmp(60644) := x"8820";
    tmp(60645) := x"8020";
    tmp(60646) := x"6800";
    tmp(60647) := x"8000";
    tmp(60648) := x"9800";
    tmp(60649) := x"a820";
    tmp(60650) := x"c020";
    tmp(60651) := x"b000";
    tmp(60652) := x"c020";
    tmp(60653) := x"a820";
    tmp(60654) := x"a000";
    tmp(60655) := x"c020";
    tmp(60656) := x"a800";
    tmp(60657) := x"b000";
    tmp(60658) := x"b800";
    tmp(60659) := x"b820";
    tmp(60660) := x"9000";
    tmp(60661) := x"a820";
    tmp(60662) := x"4861";
    tmp(60663) := x"1061";
    tmp(60664) := x"1081";
    tmp(60665) := x"1081";
    tmp(60666) := x"10a2";
    tmp(60667) := x"18a2";
    tmp(60668) := x"18c3";
    tmp(60669) := x"18e3";
    tmp(60670) := x"20e4";
    tmp(60671) := x"20e4";
    tmp(60672) := x"2104";
    tmp(60673) := x"2125";
    tmp(60674) := x"2125";
    tmp(60675) := x"2925";
    tmp(60676) := x"2925";
    tmp(60677) := x"2925";
    tmp(60678) := x"2946";
    tmp(60679) := x"2966";
    tmp(60680) := x"3167";
    tmp(60681) := x"3187";
    tmp(60682) := x"3187";
    tmp(60683) := x"3187";
    tmp(60684) := x"3187";
    tmp(60685) := x"3187";
    tmp(60686) := x"3187";
    tmp(60687) := x"3187";
    tmp(60688) := x"3187";
    tmp(60689) := x"3167";
    tmp(60690) := x"3187";
    tmp(60691) := x"3187";
    tmp(60692) := x"3187";
    tmp(60693) := x"3187";
    tmp(60694) := x"3187";
    tmp(60695) := x"3187";
    tmp(60696) := x"3187";
    tmp(60697) := x"3187";
    tmp(60698) := x"3187";
    tmp(60699) := x"3187";
    tmp(60700) := x"3187";
    tmp(60701) := x"3187";
    tmp(60702) := x"3187";
    tmp(60703) := x"3188";
    tmp(60704) := x"31a8";
    tmp(60705) := x"31a7";
    tmp(60706) := x"31a7";
    tmp(60707) := x"3187";
    tmp(60708) := x"2986";
    tmp(60709) := x"2986";
    tmp(60710) := x"2966";
    tmp(60711) := x"2965";
    tmp(60712) := x"2145";
    tmp(60713) := x"2124";
    tmp(60714) := x"2124";
    tmp(60715) := x"2124";
    tmp(60716) := x"1904";
    tmp(60717) := x"1903";
    tmp(60718) := x"1903";
    tmp(60719) := x"18e3";
    tmp(60720) := x"0000";
    tmp(60721) := x"0800";
    tmp(60722) := x"0800";
    tmp(60723) := x"0800";
    tmp(60724) := x"0800";
    tmp(60725) := x"0800";
    tmp(60726) := x"0800";
    tmp(60727) := x"0800";
    tmp(60728) := x"0800";
    tmp(60729) := x"1000";
    tmp(60730) := x"1000";
    tmp(60731) := x"1000";
    tmp(60732) := x"1000";
    tmp(60733) := x"1000";
    tmp(60734) := x"1000";
    tmp(60735) := x"1000";
    tmp(60736) := x"1000";
    tmp(60737) := x"1000";
    tmp(60738) := x"1000";
    tmp(60739) := x"1000";
    tmp(60740) := x"1000";
    tmp(60741) := x"1000";
    tmp(60742) := x"1000";
    tmp(60743) := x"1000";
    tmp(60744) := x"1000";
    tmp(60745) := x"1800";
    tmp(60746) := x"1800";
    tmp(60747) := x"1800";
    tmp(60748) := x"1800";
    tmp(60749) := x"1800";
    tmp(60750) := x"2000";
    tmp(60751) := x"2000";
    tmp(60752) := x"2000";
    tmp(60753) := x"2000";
    tmp(60754) := x"2000";
    tmp(60755) := x"2000";
    tmp(60756) := x"2000";
    tmp(60757) := x"2000";
    tmp(60758) := x"2000";
    tmp(60759) := x"2000";
    tmp(60760) := x"2000";
    tmp(60761) := x"2000";
    tmp(60762) := x"2000";
    tmp(60763) := x"2000";
    tmp(60764) := x"2000";
    tmp(60765) := x"2000";
    tmp(60766) := x"2000";
    tmp(60767) := x"2000";
    tmp(60768) := x"2000";
    tmp(60769) := x"2000";
    tmp(60770) := x"2000";
    tmp(60771) := x"2000";
    tmp(60772) := x"2000";
    tmp(60773) := x"2000";
    tmp(60774) := x"2000";
    tmp(60775) := x"2800";
    tmp(60776) := x"2800";
    tmp(60777) := x"2800";
    tmp(60778) := x"2800";
    tmp(60779) := x"2800";
    tmp(60780) := x"2800";
    tmp(60781) := x"2800";
    tmp(60782) := x"2800";
    tmp(60783) := x"3000";
    tmp(60784) := x"3000";
    tmp(60785) := x"2800";
    tmp(60786) := x"2800";
    tmp(60787) := x"2800";
    tmp(60788) := x"2800";
    tmp(60789) := x"2000";
    tmp(60790) := x"2000";
    tmp(60791) := x"1800";
    tmp(60792) := x"1000";
    tmp(60793) := x"1000";
    tmp(60794) := x"1000";
    tmp(60795) := x"1800";
    tmp(60796) := x"2000";
    tmp(60797) := x"2000";
    tmp(60798) := x"2000";
    tmp(60799) := x"1800";
    tmp(60800) := x"2000";
    tmp(60801) := x"2000";
    tmp(60802) := x"2000";
    tmp(60803) := x"2000";
    tmp(60804) := x"2000";
    tmp(60805) := x"1800";
    tmp(60806) := x"1000";
    tmp(60807) := x"1000";
    tmp(60808) := x"1000";
    tmp(60809) := x"1000";
    tmp(60810) := x"1000";
    tmp(60811) := x"1000";
    tmp(60812) := x"1000";
    tmp(60813) := x"1800";
    tmp(60814) := x"1000";
    tmp(60815) := x"1800";
    tmp(60816) := x"1800";
    tmp(60817) := x"1800";
    tmp(60818) := x"2800";
    tmp(60819) := x"2800";
    tmp(60820) := x"2800";
    tmp(60821) := x"2800";
    tmp(60822) := x"2800";
    tmp(60823) := x"2800";
    tmp(60824) := x"2800";
    tmp(60825) := x"3800";
    tmp(60826) := x"3800";
    tmp(60827) := x"4000";
    tmp(60828) := x"4800";
    tmp(60829) := x"4800";
    tmp(60830) := x"4800";
    tmp(60831) := x"5000";
    tmp(60832) := x"4800";
    tmp(60833) := x"4800";
    tmp(60834) := x"5000";
    tmp(60835) := x"5000";
    tmp(60836) := x"4800";
    tmp(60837) := x"4800";
    tmp(60838) := x"4800";
    tmp(60839) := x"4000";
    tmp(60840) := x"4000";
    tmp(60841) := x"4800";
    tmp(60842) := x"4800";
    tmp(60843) := x"5000";
    tmp(60844) := x"5000";
    tmp(60845) := x"5800";
    tmp(60846) := x"5800";
    tmp(60847) := x"5800";
    tmp(60848) := x"5800";
    tmp(60849) := x"5000";
    tmp(60850) := x"5000";
    tmp(60851) := x"6000";
    tmp(60852) := x"6800";
    tmp(60853) := x"6000";
    tmp(60854) := x"6000";
    tmp(60855) := x"6800";
    tmp(60856) := x"7000";
    tmp(60857) := x"6800";
    tmp(60858) := x"7800";
    tmp(60859) := x"8020";
    tmp(60860) := x"8820";
    tmp(60861) := x"6000";
    tmp(60862) := x"6020";
    tmp(60863) := x"6020";
    tmp(60864) := x"6820";
    tmp(60865) := x"6820";
    tmp(60866) := x"5800";
    tmp(60867) := x"6820";
    tmp(60868) := x"6020";
    tmp(60869) := x"7820";
    tmp(60870) := x"8820";
    tmp(60871) := x"6820";
    tmp(60872) := x"6820";
    tmp(60873) := x"6020";
    tmp(60874) := x"7020";
    tmp(60875) := x"7820";
    tmp(60876) := x"8820";
    tmp(60877) := x"8820";
    tmp(60878) := x"9020";
    tmp(60879) := x"8820";
    tmp(60880) := x"9020";
    tmp(60881) := x"9020";
    tmp(60882) := x"a020";
    tmp(60883) := x"9020";
    tmp(60884) := x"9020";
    tmp(60885) := x"7820";
    tmp(60886) := x"6800";
    tmp(60887) := x"7800";
    tmp(60888) := x"9000";
    tmp(60889) := x"a820";
    tmp(60890) := x"c820";
    tmp(60891) := x"b000";
    tmp(60892) := x"b820";
    tmp(60893) := x"9800";
    tmp(60894) := x"9800";
    tmp(60895) := x"b800";
    tmp(60896) := x"b000";
    tmp(60897) := x"a800";
    tmp(60898) := x"b000";
    tmp(60899) := x"a800";
    tmp(60900) := x"8800";
    tmp(60901) := x"8820";
    tmp(60902) := x"2861";
    tmp(60903) := x"1061";
    tmp(60904) := x"1081";
    tmp(60905) := x"1082";
    tmp(60906) := x"10a2";
    tmp(60907) := x"18c2";
    tmp(60908) := x"18c3";
    tmp(60909) := x"20e3";
    tmp(60910) := x"2104";
    tmp(60911) := x"2104";
    tmp(60912) := x"2104";
    tmp(60913) := x"2925";
    tmp(60914) := x"2125";
    tmp(60915) := x"2125";
    tmp(60916) := x"2925";
    tmp(60917) := x"2926";
    tmp(60918) := x"2946";
    tmp(60919) := x"2966";
    tmp(60920) := x"3167";
    tmp(60921) := x"3166";
    tmp(60922) := x"3166";
    tmp(60923) := x"3167";
    tmp(60924) := x"3167";
    tmp(60925) := x"3167";
    tmp(60926) := x"3167";
    tmp(60927) := x"3187";
    tmp(60928) := x"3187";
    tmp(60929) := x"2967";
    tmp(60930) := x"2967";
    tmp(60931) := x"2987";
    tmp(60932) := x"2967";
    tmp(60933) := x"3187";
    tmp(60934) := x"3187";
    tmp(60935) := x"3187";
    tmp(60936) := x"3187";
    tmp(60937) := x"31a7";
    tmp(60938) := x"3187";
    tmp(60939) := x"31a7";
    tmp(60940) := x"31a7";
    tmp(60941) := x"31a8";
    tmp(60942) := x"31c8";
    tmp(60943) := x"39c9";
    tmp(60944) := x"39c9";
    tmp(60945) := x"39e9";
    tmp(60946) := x"3a09";
    tmp(60947) := x"39e8";
    tmp(60948) := x"31c8";
    tmp(60949) := x"31a7";
    tmp(60950) := x"31a7";
    tmp(60951) := x"2986";
    tmp(60952) := x"2966";
    tmp(60953) := x"2965";
    tmp(60954) := x"2965";
    tmp(60955) := x"2145";
    tmp(60956) := x"2145";
    tmp(60957) := x"2144";
    tmp(60958) := x"2124";
    tmp(60959) := x"1923";
    tmp(60960) := x"0000";
    tmp(60961) := x"0800";
    tmp(60962) := x"0800";
    tmp(60963) := x"0800";
    tmp(60964) := x"0800";
    tmp(60965) := x"0800";
    tmp(60966) := x"0800";
    tmp(60967) := x"0800";
    tmp(60968) := x"0800";
    tmp(60969) := x"1000";
    tmp(60970) := x"1000";
    tmp(60971) := x"1000";
    tmp(60972) := x"1000";
    tmp(60973) := x"1000";
    tmp(60974) := x"1000";
    tmp(60975) := x"1000";
    tmp(60976) := x"1000";
    tmp(60977) := x"1000";
    tmp(60978) := x"1000";
    tmp(60979) := x"1000";
    tmp(60980) := x"1000";
    tmp(60981) := x"1000";
    tmp(60982) := x"1800";
    tmp(60983) := x"1800";
    tmp(60984) := x"1800";
    tmp(60985) := x"1800";
    tmp(60986) := x"1800";
    tmp(60987) := x"1800";
    tmp(60988) := x"1800";
    tmp(60989) := x"2000";
    tmp(60990) := x"2000";
    tmp(60991) := x"2000";
    tmp(60992) := x"2000";
    tmp(60993) := x"2000";
    tmp(60994) := x"2000";
    tmp(60995) := x"2000";
    tmp(60996) := x"1800";
    tmp(60997) := x"1800";
    tmp(60998) := x"2000";
    tmp(60999) := x"1800";
    tmp(61000) := x"2000";
    tmp(61001) := x"2000";
    tmp(61002) := x"2000";
    tmp(61003) := x"2000";
    tmp(61004) := x"2000";
    tmp(61005) := x"2000";
    tmp(61006) := x"2800";
    tmp(61007) := x"2000";
    tmp(61008) := x"2000";
    tmp(61009) := x"2000";
    tmp(61010) := x"2000";
    tmp(61011) := x"2800";
    tmp(61012) := x"2800";
    tmp(61013) := x"2800";
    tmp(61014) := x"2800";
    tmp(61015) := x"2800";
    tmp(61016) := x"2800";
    tmp(61017) := x"3000";
    tmp(61018) := x"2800";
    tmp(61019) := x"2800";
    tmp(61020) := x"2800";
    tmp(61021) := x"2800";
    tmp(61022) := x"2800";
    tmp(61023) := x"2800";
    tmp(61024) := x"3000";
    tmp(61025) := x"3000";
    tmp(61026) := x"2800";
    tmp(61027) := x"2800";
    tmp(61028) := x"2800";
    tmp(61029) := x"2800";
    tmp(61030) := x"2000";
    tmp(61031) := x"1000";
    tmp(61032) := x"0800";
    tmp(61033) := x"1000";
    tmp(61034) := x"1000";
    tmp(61035) := x"1000";
    tmp(61036) := x"1800";
    tmp(61037) := x"1800";
    tmp(61038) := x"1800";
    tmp(61039) := x"2000";
    tmp(61040) := x"2000";
    tmp(61041) := x"2000";
    tmp(61042) := x"2000";
    tmp(61043) := x"2000";
    tmp(61044) := x"2000";
    tmp(61045) := x"1800";
    tmp(61046) := x"1000";
    tmp(61047) := x"1000";
    tmp(61048) := x"1000";
    tmp(61049) := x"1000";
    tmp(61050) := x"1000";
    tmp(61051) := x"1000";
    tmp(61052) := x"1800";
    tmp(61053) := x"1800";
    tmp(61054) := x"1800";
    tmp(61055) := x"1800";
    tmp(61056) := x"1800";
    tmp(61057) := x"2000";
    tmp(61058) := x"2000";
    tmp(61059) := x"2000";
    tmp(61060) := x"2000";
    tmp(61061) := x"1800";
    tmp(61062) := x"1800";
    tmp(61063) := x"1800";
    tmp(61064) := x"2000";
    tmp(61065) := x"2800";
    tmp(61066) := x"2800";
    tmp(61067) := x"3800";
    tmp(61068) := x"4000";
    tmp(61069) := x"4800";
    tmp(61070) := x"5000";
    tmp(61071) := x"5000";
    tmp(61072) := x"4800";
    tmp(61073) := x"4800";
    tmp(61074) := x"5000";
    tmp(61075) := x"5000";
    tmp(61076) := x"5000";
    tmp(61077) := x"5000";
    tmp(61078) := x"4800";
    tmp(61079) := x"4000";
    tmp(61080) := x"4800";
    tmp(61081) := x"4800";
    tmp(61082) := x"4800";
    tmp(61083) := x"5000";
    tmp(61084) := x"5000";
    tmp(61085) := x"5000";
    tmp(61086) := x"5800";
    tmp(61087) := x"5800";
    tmp(61088) := x"5000";
    tmp(61089) := x"5800";
    tmp(61090) := x"5800";
    tmp(61091) := x"6000";
    tmp(61092) := x"6800";
    tmp(61093) := x"5800";
    tmp(61094) := x"6000";
    tmp(61095) := x"6800";
    tmp(61096) := x"6800";
    tmp(61097) := x"7000";
    tmp(61098) := x"7800";
    tmp(61099) := x"8020";
    tmp(61100) := x"9020";
    tmp(61101) := x"6000";
    tmp(61102) := x"6000";
    tmp(61103) := x"6820";
    tmp(61104) := x"6820";
    tmp(61105) := x"6820";
    tmp(61106) := x"5820";
    tmp(61107) := x"6820";
    tmp(61108) := x"6000";
    tmp(61109) := x"6820";
    tmp(61110) := x"9040";
    tmp(61111) := x"7020";
    tmp(61112) := x"7020";
    tmp(61113) := x"6820";
    tmp(61114) := x"6820";
    tmp(61115) := x"7820";
    tmp(61116) := x"8820";
    tmp(61117) := x"8820";
    tmp(61118) := x"8820";
    tmp(61119) := x"8820";
    tmp(61120) := x"a040";
    tmp(61121) := x"9840";
    tmp(61122) := x"a020";
    tmp(61123) := x"9020";
    tmp(61124) := x"8820";
    tmp(61125) := x"8020";
    tmp(61126) := x"6800";
    tmp(61127) := x"7000";
    tmp(61128) := x"8800";
    tmp(61129) := x"9820";
    tmp(61130) := x"b820";
    tmp(61131) := x"b820";
    tmp(61132) := x"b000";
    tmp(61133) := x"9000";
    tmp(61134) := x"9000";
    tmp(61135) := x"b000";
    tmp(61136) := x"a000";
    tmp(61137) := x"9800";
    tmp(61138) := x"b820";
    tmp(61139) := x"a000";
    tmp(61140) := x"9000";
    tmp(61141) := x"7040";
    tmp(61142) := x"1861";
    tmp(61143) := x"1061";
    tmp(61144) := x"1081";
    tmp(61145) := x"1082";
    tmp(61146) := x"18a2";
    tmp(61147) := x"18c3";
    tmp(61148) := x"18e3";
    tmp(61149) := x"20e4";
    tmp(61150) := x"2104";
    tmp(61151) := x"2104";
    tmp(61152) := x"2104";
    tmp(61153) := x"2105";
    tmp(61154) := x"2125";
    tmp(61155) := x"2125";
    tmp(61156) := x"2925";
    tmp(61157) := x"2925";
    tmp(61158) := x"2946";
    tmp(61159) := x"2966";
    tmp(61160) := x"2966";
    tmp(61161) := x"2966";
    tmp(61162) := x"2966";
    tmp(61163) := x"2966";
    tmp(61164) := x"2946";
    tmp(61165) := x"2966";
    tmp(61166) := x"2966";
    tmp(61167) := x"2966";
    tmp(61168) := x"2967";
    tmp(61169) := x"2966";
    tmp(61170) := x"2966";
    tmp(61171) := x"2967";
    tmp(61172) := x"3167";
    tmp(61173) := x"3187";
    tmp(61174) := x"3187";
    tmp(61175) := x"3187";
    tmp(61176) := x"31a8";
    tmp(61177) := x"31a8";
    tmp(61178) := x"31a8";
    tmp(61179) := x"31a8";
    tmp(61180) := x"31a8";
    tmp(61181) := x"39e9";
    tmp(61182) := x"39ea";
    tmp(61183) := x"3a0a";
    tmp(61184) := x"424b";
    tmp(61185) := x"422a";
    tmp(61186) := x"422a";
    tmp(61187) := x"422a";
    tmp(61188) := x"3a09";
    tmp(61189) := x"39e9";
    tmp(61190) := x"39e8";
    tmp(61191) := x"31e8";
    tmp(61192) := x"31a7";
    tmp(61193) := x"31a6";
    tmp(61194) := x"31a6";
    tmp(61195) := x"2986";
    tmp(61196) := x"2985";
    tmp(61197) := x"2965";
    tmp(61198) := x"2165";
    tmp(61199) := x"2164";
    tmp(61200) := x"0000";
    tmp(61201) := x"0800";
    tmp(61202) := x"0800";
    tmp(61203) := x"0800";
    tmp(61204) := x"0800";
    tmp(61205) := x"0800";
    tmp(61206) := x"0800";
    tmp(61207) := x"0800";
    tmp(61208) := x"0800";
    tmp(61209) := x"0800";
    tmp(61210) := x"1000";
    tmp(61211) := x"1000";
    tmp(61212) := x"1000";
    tmp(61213) := x"1000";
    tmp(61214) := x"1000";
    tmp(61215) := x"1000";
    tmp(61216) := x"1000";
    tmp(61217) := x"1000";
    tmp(61218) := x"1000";
    tmp(61219) := x"1000";
    tmp(61220) := x"1000";
    tmp(61221) := x"1000";
    tmp(61222) := x"1800";
    tmp(61223) := x"1800";
    tmp(61224) := x"1800";
    tmp(61225) := x"1800";
    tmp(61226) := x"1800";
    tmp(61227) := x"1800";
    tmp(61228) := x"2000";
    tmp(61229) := x"2000";
    tmp(61230) := x"2000";
    tmp(61231) := x"2000";
    tmp(61232) := x"2000";
    tmp(61233) := x"2000";
    tmp(61234) := x"2000";
    tmp(61235) := x"2000";
    tmp(61236) := x"1800";
    tmp(61237) := x"1800";
    tmp(61238) := x"1800";
    tmp(61239) := x"1800";
    tmp(61240) := x"1800";
    tmp(61241) := x"2000";
    tmp(61242) := x"2000";
    tmp(61243) := x"2000";
    tmp(61244) := x"2800";
    tmp(61245) := x"2800";
    tmp(61246) := x"2800";
    tmp(61247) := x"2800";
    tmp(61248) := x"2000";
    tmp(61249) := x"2000";
    tmp(61250) := x"2000";
    tmp(61251) := x"2800";
    tmp(61252) := x"2800";
    tmp(61253) := x"2800";
    tmp(61254) := x"2800";
    tmp(61255) := x"3000";
    tmp(61256) := x"3000";
    tmp(61257) := x"3000";
    tmp(61258) := x"3000";
    tmp(61259) := x"2800";
    tmp(61260) := x"2800";
    tmp(61261) := x"3000";
    tmp(61262) := x"3000";
    tmp(61263) := x"2800";
    tmp(61264) := x"3000";
    tmp(61265) := x"3000";
    tmp(61266) := x"3000";
    tmp(61267) := x"2800";
    tmp(61268) := x"2800";
    tmp(61269) := x"2000";
    tmp(61270) := x"1000";
    tmp(61271) := x"0800";
    tmp(61272) := x"0800";
    tmp(61273) := x"0800";
    tmp(61274) := x"0800";
    tmp(61275) := x"1000";
    tmp(61276) := x"1000";
    tmp(61277) := x"1000";
    tmp(61278) := x"1800";
    tmp(61279) := x"1800";
    tmp(61280) := x"1800";
    tmp(61281) := x"2000";
    tmp(61282) := x"2000";
    tmp(61283) := x"1800";
    tmp(61284) := x"1800";
    tmp(61285) := x"1800";
    tmp(61286) := x"1000";
    tmp(61287) := x"1000";
    tmp(61288) := x"1000";
    tmp(61289) := x"1000";
    tmp(61290) := x"1000";
    tmp(61291) := x"1000";
    tmp(61292) := x"1800";
    tmp(61293) := x"1800";
    tmp(61294) := x"1800";
    tmp(61295) := x"1800";
    tmp(61296) := x"1800";
    tmp(61297) := x"1800";
    tmp(61298) := x"1800";
    tmp(61299) := x"1800";
    tmp(61300) := x"1000";
    tmp(61301) := x"1000";
    tmp(61302) := x"1000";
    tmp(61303) := x"1800";
    tmp(61304) := x"2000";
    tmp(61305) := x"2800";
    tmp(61306) := x"2800";
    tmp(61307) := x"3000";
    tmp(61308) := x"3800";
    tmp(61309) := x"4000";
    tmp(61310) := x"4000";
    tmp(61311) := x"4800";
    tmp(61312) := x"4800";
    tmp(61313) := x"5000";
    tmp(61314) := x"4800";
    tmp(61315) := x"4800";
    tmp(61316) := x"5000";
    tmp(61317) := x"5000";
    tmp(61318) := x"4800";
    tmp(61319) := x"4000";
    tmp(61320) := x"4000";
    tmp(61321) := x"4000";
    tmp(61322) := x"4800";
    tmp(61323) := x"5000";
    tmp(61324) := x"4800";
    tmp(61325) := x"5000";
    tmp(61326) := x"5000";
    tmp(61327) := x"5800";
    tmp(61328) := x"5800";
    tmp(61329) := x"5800";
    tmp(61330) := x"5800";
    tmp(61331) := x"6800";
    tmp(61332) := x"6000";
    tmp(61333) := x"5800";
    tmp(61334) := x"6000";
    tmp(61335) := x"6800";
    tmp(61336) := x"6800";
    tmp(61337) := x"7000";
    tmp(61338) := x"7000";
    tmp(61339) := x"8020";
    tmp(61340) := x"9020";
    tmp(61341) := x"6800";
    tmp(61342) := x"6000";
    tmp(61343) := x"6820";
    tmp(61344) := x"6820";
    tmp(61345) := x"6820";
    tmp(61346) := x"5820";
    tmp(61347) := x"6820";
    tmp(61348) := x"6820";
    tmp(61349) := x"6820";
    tmp(61350) := x"8020";
    tmp(61351) := x"7820";
    tmp(61352) := x"7820";
    tmp(61353) := x"6020";
    tmp(61354) := x"6020";
    tmp(61355) := x"8020";
    tmp(61356) := x"8820";
    tmp(61357) := x"8820";
    tmp(61358) := x"8820";
    tmp(61359) := x"9020";
    tmp(61360) := x"9020";
    tmp(61361) := x"a040";
    tmp(61362) := x"8820";
    tmp(61363) := x"9020";
    tmp(61364) := x"8820";
    tmp(61365) := x"7820";
    tmp(61366) := x"6800";
    tmp(61367) := x"7000";
    tmp(61368) := x"8000";
    tmp(61369) := x"9000";
    tmp(61370) := x"b020";
    tmp(61371) := x"b820";
    tmp(61372) := x"a820";
    tmp(61373) := x"9000";
    tmp(61374) := x"8800";
    tmp(61375) := x"a800";
    tmp(61376) := x"a000";
    tmp(61377) := x"9800";
    tmp(61378) := x"b820";
    tmp(61379) := x"9000";
    tmp(61380) := x"9020";
    tmp(61381) := x"3841";
    tmp(61382) := x"1061";
    tmp(61383) := x"1081";
    tmp(61384) := x"1082";
    tmp(61385) := x"10a2";
    tmp(61386) := x"18a2";
    tmp(61387) := x"18c3";
    tmp(61388) := x"18e3";
    tmp(61389) := x"20e4";
    tmp(61390) := x"2104";
    tmp(61391) := x"2104";
    tmp(61392) := x"2104";
    tmp(61393) := x"2105";
    tmp(61394) := x"2104";
    tmp(61395) := x"2104";
    tmp(61396) := x"2125";
    tmp(61397) := x"2925";
    tmp(61398) := x"2925";
    tmp(61399) := x"2926";
    tmp(61400) := x"2926";
    tmp(61401) := x"2946";
    tmp(61402) := x"2946";
    tmp(61403) := x"2946";
    tmp(61404) := x"2926";
    tmp(61405) := x"2946";
    tmp(61406) := x"2946";
    tmp(61407) := x"2966";
    tmp(61408) := x"2966";
    tmp(61409) := x"2966";
    tmp(61410) := x"2966";
    tmp(61411) := x"3187";
    tmp(61412) := x"3187";
    tmp(61413) := x"3187";
    tmp(61414) := x"3187";
    tmp(61415) := x"31a7";
    tmp(61416) := x"31a8";
    tmp(61417) := x"39c8";
    tmp(61418) := x"39c8";
    tmp(61419) := x"39c8";
    tmp(61420) := x"39e9";
    tmp(61421) := x"4209";
    tmp(61422) := x"422a";
    tmp(61423) := x"422b";
    tmp(61424) := x"424b";
    tmp(61425) := x"424b";
    tmp(61426) := x"4a6b";
    tmp(61427) := x"4a6b";
    tmp(61428) := x"4a6b";
    tmp(61429) := x"424a";
    tmp(61430) := x"3a29";
    tmp(61431) := x"3a09";
    tmp(61432) := x"39e8";
    tmp(61433) := x"31c7";
    tmp(61434) := x"31c7";
    tmp(61435) := x"31a6";
    tmp(61436) := x"31a6";
    tmp(61437) := x"2986";
    tmp(61438) := x"2985";
    tmp(61439) := x"2985";
    tmp(61440) := x"0000";
    tmp(61441) := x"0800";
    tmp(61442) := x"0800";
    tmp(61443) := x"0800";
    tmp(61444) := x"0800";
    tmp(61445) := x"0800";
    tmp(61446) := x"0800";
    tmp(61447) := x"0800";
    tmp(61448) := x"0800";
    tmp(61449) := x"1000";
    tmp(61450) := x"1000";
    tmp(61451) := x"1000";
    tmp(61452) := x"1000";
    tmp(61453) := x"1000";
    tmp(61454) := x"1000";
    tmp(61455) := x"1000";
    tmp(61456) := x"1000";
    tmp(61457) := x"1000";
    tmp(61458) := x"1000";
    tmp(61459) := x"1000";
    tmp(61460) := x"1000";
    tmp(61461) := x"1000";
    tmp(61462) := x"1000";
    tmp(61463) := x"1800";
    tmp(61464) := x"1800";
    tmp(61465) := x"1800";
    tmp(61466) := x"1800";
    tmp(61467) := x"1800";
    tmp(61468) := x"1800";
    tmp(61469) := x"1800";
    tmp(61470) := x"2000";
    tmp(61471) := x"2000";
    tmp(61472) := x"2800";
    tmp(61473) := x"2000";
    tmp(61474) := x"2000";
    tmp(61475) := x"1800";
    tmp(61476) := x"1800";
    tmp(61477) := x"1800";
    tmp(61478) := x"1800";
    tmp(61479) := x"1800";
    tmp(61480) := x"1800";
    tmp(61481) := x"2000";
    tmp(61482) := x"2000";
    tmp(61483) := x"2000";
    tmp(61484) := x"2000";
    tmp(61485) := x"2800";
    tmp(61486) := x"2800";
    tmp(61487) := x"2800";
    tmp(61488) := x"2000";
    tmp(61489) := x"2000";
    tmp(61490) := x"2000";
    tmp(61491) := x"2000";
    tmp(61492) := x"2800";
    tmp(61493) := x"2800";
    tmp(61494) := x"2800";
    tmp(61495) := x"2800";
    tmp(61496) := x"2800";
    tmp(61497) := x"3000";
    tmp(61498) := x"2800";
    tmp(61499) := x"2800";
    tmp(61500) := x"3000";
    tmp(61501) := x"3000";
    tmp(61502) := x"3000";
    tmp(61503) := x"3000";
    tmp(61504) := x"3000";
    tmp(61505) := x"3000";
    tmp(61506) := x"3000";
    tmp(61507) := x"2800";
    tmp(61508) := x"1820";
    tmp(61509) := x"1020";
    tmp(61510) := x"1000";
    tmp(61511) := x"0800";
    tmp(61512) := x"0800";
    tmp(61513) := x"0800";
    tmp(61514) := x"0800";
    tmp(61515) := x"0800";
    tmp(61516) := x"0800";
    tmp(61517) := x"0800";
    tmp(61518) := x"1000";
    tmp(61519) := x"1000";
    tmp(61520) := x"1000";
    tmp(61521) := x"1800";
    tmp(61522) := x"1800";
    tmp(61523) := x"1800";
    tmp(61524) := x"1800";
    tmp(61525) := x"1000";
    tmp(61526) := x"1000";
    tmp(61527) := x"1000";
    tmp(61528) := x"1000";
    tmp(61529) := x"1000";
    tmp(61530) := x"1000";
    tmp(61531) := x"1000";
    tmp(61532) := x"1000";
    tmp(61533) := x"1800";
    tmp(61534) := x"2000";
    tmp(61535) := x"2000";
    tmp(61536) := x"2000";
    tmp(61537) := x"1800";
    tmp(61538) := x"1800";
    tmp(61539) := x"1800";
    tmp(61540) := x"1000";
    tmp(61541) := x"1000";
    tmp(61542) := x"1800";
    tmp(61543) := x"2000";
    tmp(61544) := x"2800";
    tmp(61545) := x"2000";
    tmp(61546) := x"2000";
    tmp(61547) := x"2800";
    tmp(61548) := x"2800";
    tmp(61549) := x"4000";
    tmp(61550) := x"4000";
    tmp(61551) := x"4800";
    tmp(61552) := x"5000";
    tmp(61553) := x"5000";
    tmp(61554) := x"5000";
    tmp(61555) := x"5000";
    tmp(61556) := x"4800";
    tmp(61557) := x"5000";
    tmp(61558) := x"4800";
    tmp(61559) := x"4000";
    tmp(61560) := x"4000";
    tmp(61561) := x"4000";
    tmp(61562) := x"4800";
    tmp(61563) := x"4800";
    tmp(61564) := x"4800";
    tmp(61565) := x"5000";
    tmp(61566) := x"5000";
    tmp(61567) := x"5800";
    tmp(61568) := x"6000";
    tmp(61569) := x"6000";
    tmp(61570) := x"6000";
    tmp(61571) := x"6000";
    tmp(61572) := x"6000";
    tmp(61573) := x"6000";
    tmp(61574) := x"6000";
    tmp(61575) := x"6000";
    tmp(61576) := x"6800";
    tmp(61577) := x"6800";
    tmp(61578) := x"7800";
    tmp(61579) := x"8020";
    tmp(61580) := x"8820";
    tmp(61581) := x"6000";
    tmp(61582) := x"5800";
    tmp(61583) := x"6820";
    tmp(61584) := x"7020";
    tmp(61585) := x"6020";
    tmp(61586) := x"6020";
    tmp(61587) := x"6820";
    tmp(61588) := x"6820";
    tmp(61589) := x"6820";
    tmp(61590) := x"7820";
    tmp(61591) := x"8820";
    tmp(61592) := x"7020";
    tmp(61593) := x"6820";
    tmp(61594) := x"6020";
    tmp(61595) := x"8020";
    tmp(61596) := x"8820";
    tmp(61597) := x"8820";
    tmp(61598) := x"8820";
    tmp(61599) := x"9820";
    tmp(61600) := x"8820";
    tmp(61601) := x"a040";
    tmp(61602) := x"8820";
    tmp(61603) := x"9820";
    tmp(61604) := x"9020";
    tmp(61605) := x"8020";
    tmp(61606) := x"7000";
    tmp(61607) := x"7000";
    tmp(61608) := x"8000";
    tmp(61609) := x"9000";
    tmp(61610) := x"a820";
    tmp(61611) := x"b820";
    tmp(61612) := x"a820";
    tmp(61613) := x"9000";
    tmp(61614) := x"9000";
    tmp(61615) := x"a800";
    tmp(61616) := x"a000";
    tmp(61617) := x"9800";
    tmp(61618) := x"c020";
    tmp(61619) := x"9800";
    tmp(61620) := x"7020";
    tmp(61621) := x"2041";
    tmp(61622) := x"1061";
    tmp(61623) := x"1081";
    tmp(61624) := x"1082";
    tmp(61625) := x"18a2";
    tmp(61626) := x"18c2";
    tmp(61627) := x"18c3";
    tmp(61628) := x"18e3";
    tmp(61629) := x"18e4";
    tmp(61630) := x"18e4";
    tmp(61631) := x"20e4";
    tmp(61632) := x"20e4";
    tmp(61633) := x"20e4";
    tmp(61634) := x"20e4";
    tmp(61635) := x"2104";
    tmp(61636) := x"2104";
    tmp(61637) := x"2105";
    tmp(61638) := x"2925";
    tmp(61639) := x"2125";
    tmp(61640) := x"2125";
    tmp(61641) := x"2925";
    tmp(61642) := x"2925";
    tmp(61643) := x"2925";
    tmp(61644) := x"2925";
    tmp(61645) := x"2945";
    tmp(61646) := x"2925";
    tmp(61647) := x"2946";
    tmp(61648) := x"2966";
    tmp(61649) := x"2966";
    tmp(61650) := x"3167";
    tmp(61651) := x"3187";
    tmp(61652) := x"3167";
    tmp(61653) := x"3187";
    tmp(61654) := x"31a7";
    tmp(61655) := x"31a7";
    tmp(61656) := x"39c8";
    tmp(61657) := x"39e9";
    tmp(61658) := x"39e9";
    tmp(61659) := x"41e9";
    tmp(61660) := x"422a";
    tmp(61661) := x"422a";
    tmp(61662) := x"422a";
    tmp(61663) := x"4a2b";
    tmp(61664) := x"4a4b";
    tmp(61665) := x"4a4b";
    tmp(61666) := x"4a6b";
    tmp(61667) := x"4a6b";
    tmp(61668) := x"4a6b";
    tmp(61669) := x"424a";
    tmp(61670) := x"4229";
    tmp(61671) := x"3a29";
    tmp(61672) := x"3a08";
    tmp(61673) := x"39e8";
    tmp(61674) := x"39e8";
    tmp(61675) := x"39e7";
    tmp(61676) := x"31e7";
    tmp(61677) := x"31c7";
    tmp(61678) := x"31c6";
    tmp(61679) := x"29a6";
    tmp(61680) := x"0000";
    tmp(61681) := x"0800";
    tmp(61682) := x"0800";
    tmp(61683) := x"0800";
    tmp(61684) := x"0800";
    tmp(61685) := x"0800";
    tmp(61686) := x"0800";
    tmp(61687) := x"0800";
    tmp(61688) := x"1000";
    tmp(61689) := x"1000";
    tmp(61690) := x"1000";
    tmp(61691) := x"1000";
    tmp(61692) := x"1000";
    tmp(61693) := x"1000";
    tmp(61694) := x"1000";
    tmp(61695) := x"1000";
    tmp(61696) := x"1000";
    tmp(61697) := x"1000";
    tmp(61698) := x"1000";
    tmp(61699) := x"1000";
    tmp(61700) := x"1000";
    tmp(61701) := x"1000";
    tmp(61702) := x"1000";
    tmp(61703) := x"1800";
    tmp(61704) := x"1800";
    tmp(61705) := x"1800";
    tmp(61706) := x"1800";
    tmp(61707) := x"1800";
    tmp(61708) := x"1800";
    tmp(61709) := x"1800";
    tmp(61710) := x"1800";
    tmp(61711) := x"1800";
    tmp(61712) := x"2000";
    tmp(61713) := x"2000";
    tmp(61714) := x"1800";
    tmp(61715) := x"1800";
    tmp(61716) := x"1800";
    tmp(61717) := x"1800";
    tmp(61718) := x"1800";
    tmp(61719) := x"1800";
    tmp(61720) := x"1800";
    tmp(61721) := x"2000";
    tmp(61722) := x"2000";
    tmp(61723) := x"2000";
    tmp(61724) := x"2000";
    tmp(61725) := x"2000";
    tmp(61726) := x"2800";
    tmp(61727) := x"2800";
    tmp(61728) := x"2000";
    tmp(61729) := x"2000";
    tmp(61730) := x"2000";
    tmp(61731) := x"2000";
    tmp(61732) := x"2000";
    tmp(61733) := x"2000";
    tmp(61734) := x"2000";
    tmp(61735) := x"2000";
    tmp(61736) := x"2800";
    tmp(61737) := x"3000";
    tmp(61738) := x"3000";
    tmp(61739) := x"3000";
    tmp(61740) := x"2800";
    tmp(61741) := x"2800";
    tmp(61742) := x"3000";
    tmp(61743) := x"3000";
    tmp(61744) := x"3000";
    tmp(61745) := x"3000";
    tmp(61746) := x"2820";
    tmp(61747) := x"2020";
    tmp(61748) := x"1820";
    tmp(61749) := x"1020";
    tmp(61750) := x"1000";
    tmp(61751) := x"0800";
    tmp(61752) := x"0800";
    tmp(61753) := x"0800";
    tmp(61754) := x"1000";
    tmp(61755) := x"1000";
    tmp(61756) := x"1020";
    tmp(61757) := x"0800";
    tmp(61758) := x"0800";
    tmp(61759) := x"0800";
    tmp(61760) := x"1000";
    tmp(61761) := x"1000";
    tmp(61762) := x"1000";
    tmp(61763) := x"1000";
    tmp(61764) := x"1000";
    tmp(61765) := x"1000";
    tmp(61766) := x"1000";
    tmp(61767) := x"1000";
    tmp(61768) := x"1000";
    tmp(61769) := x"1000";
    tmp(61770) := x"1800";
    tmp(61771) := x"1800";
    tmp(61772) := x"1800";
    tmp(61773) := x"1800";
    tmp(61774) := x"2000";
    tmp(61775) := x"2000";
    tmp(61776) := x"2000";
    tmp(61777) := x"2000";
    tmp(61778) := x"2000";
    tmp(61779) := x"2000";
    tmp(61780) := x"2000";
    tmp(61781) := x"2000";
    tmp(61782) := x"2000";
    tmp(61783) := x"1800";
    tmp(61784) := x"1800";
    tmp(61785) := x"1800";
    tmp(61786) := x"1000";
    tmp(61787) := x"1000";
    tmp(61788) := x"1800";
    tmp(61789) := x"3800";
    tmp(61790) := x"4000";
    tmp(61791) := x"4800";
    tmp(61792) := x"4800";
    tmp(61793) := x"4800";
    tmp(61794) := x"4800";
    tmp(61795) := x"5000";
    tmp(61796) := x"4800";
    tmp(61797) := x"4800";
    tmp(61798) := x"4000";
    tmp(61799) := x"4000";
    tmp(61800) := x"4000";
    tmp(61801) := x"4800";
    tmp(61802) := x"5000";
    tmp(61803) := x"4800";
    tmp(61804) := x"4800";
    tmp(61805) := x"5000";
    tmp(61806) := x"5800";
    tmp(61807) := x"5800";
    tmp(61808) := x"5800";
    tmp(61809) := x"6800";
    tmp(61810) := x"6000";
    tmp(61811) := x"5800";
    tmp(61812) := x"5800";
    tmp(61813) := x"6800";
    tmp(61814) := x"6000";
    tmp(61815) := x"6800";
    tmp(61816) := x"6000";
    tmp(61817) := x"6000";
    tmp(61818) := x"7000";
    tmp(61819) := x"8820";
    tmp(61820) := x"7020";
    tmp(61821) := x"6000";
    tmp(61822) := x"5800";
    tmp(61823) := x"6820";
    tmp(61824) := x"6820";
    tmp(61825) := x"6020";
    tmp(61826) := x"6020";
    tmp(61827) := x"7020";
    tmp(61828) := x"6820";
    tmp(61829) := x"6820";
    tmp(61830) := x"7820";
    tmp(61831) := x"9020";
    tmp(61832) := x"7020";
    tmp(61833) := x"6820";
    tmp(61834) := x"6020";
    tmp(61835) := x"7820";
    tmp(61836) := x"8820";
    tmp(61837) := x"9020";
    tmp(61838) := x"9020";
    tmp(61839) := x"9820";
    tmp(61840) := x"9020";
    tmp(61841) := x"a040";
    tmp(61842) := x"8820";
    tmp(61843) := x"9020";
    tmp(61844) := x"9020";
    tmp(61845) := x"9020";
    tmp(61846) := x"7800";
    tmp(61847) := x"7800";
    tmp(61848) := x"7800";
    tmp(61849) := x"8800";
    tmp(61850) := x"9820";
    tmp(61851) := x"a820";
    tmp(61852) := x"a020";
    tmp(61853) := x"8800";
    tmp(61854) := x"9800";
    tmp(61855) := x"a000";
    tmp(61856) := x"b020";
    tmp(61857) := x"a820";
    tmp(61858) := x"d820";
    tmp(61859) := x"9800";
    tmp(61860) := x"5020";
    tmp(61861) := x"1841";
    tmp(61862) := x"1061";
    tmp(61863) := x"1081";
    tmp(61864) := x"10a2";
    tmp(61865) := x"10a2";
    tmp(61866) := x"18a2";
    tmp(61867) := x"18c3";
    tmp(61868) := x"18c3";
    tmp(61869) := x"18c3";
    tmp(61870) := x"18c3";
    tmp(61871) := x"18c3";
    tmp(61872) := x"18c3";
    tmp(61873) := x"18e3";
    tmp(61874) := x"18e3";
    tmp(61875) := x"20e4";
    tmp(61876) := x"2104";
    tmp(61877) := x"2104";
    tmp(61878) := x"2104";
    tmp(61879) := x"2104";
    tmp(61880) := x"2104";
    tmp(61881) := x"2105";
    tmp(61882) := x"2105";
    tmp(61883) := x"2125";
    tmp(61884) := x"2925";
    tmp(61885) := x"2925";
    tmp(61886) := x"2925";
    tmp(61887) := x"2946";
    tmp(61888) := x"2946";
    tmp(61889) := x"2966";
    tmp(61890) := x"3167";
    tmp(61891) := x"3187";
    tmp(61892) := x"3187";
    tmp(61893) := x"3187";
    tmp(61894) := x"31a7";
    tmp(61895) := x"39a8";
    tmp(61896) := x"39e8";
    tmp(61897) := x"39e9";
    tmp(61898) := x"39e9";
    tmp(61899) := x"41e9";
    tmp(61900) := x"4209";
    tmp(61901) := x"422a";
    tmp(61902) := x"422a";
    tmp(61903) := x"4a4b";
    tmp(61904) := x"4a4b";
    tmp(61905) := x"4a4b";
    tmp(61906) := x"4a4b";
    tmp(61907) := x"4a6b";
    tmp(61908) := x"4a6b";
    tmp(61909) := x"4a6b";
    tmp(61910) := x"424a";
    tmp(61911) := x"4229";
    tmp(61912) := x"4229";
    tmp(61913) := x"4229";
    tmp(61914) := x"3a09";
    tmp(61915) := x"4209";
    tmp(61916) := x"4229";
    tmp(61917) := x"3a08";
    tmp(61918) := x"39e7";
    tmp(61919) := x"31e7";
    tmp(61920) := x"0000";
    tmp(61921) := x"0800";
    tmp(61922) := x"0800";
    tmp(61923) := x"0800";
    tmp(61924) := x"0800";
    tmp(61925) := x"0800";
    tmp(61926) := x"0800";
    tmp(61927) := x"0800";
    tmp(61928) := x"1000";
    tmp(61929) := x"1000";
    tmp(61930) := x"1000";
    tmp(61931) := x"1000";
    tmp(61932) := x"1000";
    tmp(61933) := x"1000";
    tmp(61934) := x"1000";
    tmp(61935) := x"1000";
    tmp(61936) := x"1000";
    tmp(61937) := x"1000";
    tmp(61938) := x"1000";
    tmp(61939) := x"1000";
    tmp(61940) := x"1000";
    tmp(61941) := x"1000";
    tmp(61942) := x"1000";
    tmp(61943) := x"1800";
    tmp(61944) := x"1800";
    tmp(61945) := x"1800";
    tmp(61946) := x"1800";
    tmp(61947) := x"1800";
    tmp(61948) := x"1800";
    tmp(61949) := x"1800";
    tmp(61950) := x"1800";
    tmp(61951) := x"1800";
    tmp(61952) := x"1800";
    tmp(61953) := x"1800";
    tmp(61954) := x"1800";
    tmp(61955) := x"1800";
    tmp(61956) := x"1800";
    tmp(61957) := x"1800";
    tmp(61958) := x"1800";
    tmp(61959) := x"1800";
    tmp(61960) := x"1800";
    tmp(61961) := x"1800";
    tmp(61962) := x"2000";
    tmp(61963) := x"2000";
    tmp(61964) := x"2000";
    tmp(61965) := x"2000";
    tmp(61966) := x"2800";
    tmp(61967) := x"2800";
    tmp(61968) := x"2000";
    tmp(61969) := x"2000";
    tmp(61970) := x"2000";
    tmp(61971) := x"2000";
    tmp(61972) := x"2000";
    tmp(61973) := x"2000";
    tmp(61974) := x"2000";
    tmp(61975) := x"2800";
    tmp(61976) := x"3000";
    tmp(61977) := x"2800";
    tmp(61978) := x"2800";
    tmp(61979) := x"3000";
    tmp(61980) := x"3000";
    tmp(61981) := x"3000";
    tmp(61982) := x"3000";
    tmp(61983) := x"3000";
    tmp(61984) := x"3000";
    tmp(61985) := x"3020";
    tmp(61986) := x"2820";
    tmp(61987) := x"2020";
    tmp(61988) := x"1800";
    tmp(61989) := x"1000";
    tmp(61990) := x"1000";
    tmp(61991) := x"1000";
    tmp(61992) := x"1800";
    tmp(61993) := x"1800";
    tmp(61994) := x"1800";
    tmp(61995) := x"1000";
    tmp(61996) := x"0800";
    tmp(61997) := x"0820";
    tmp(61998) := x"0820";
    tmp(61999) := x"0800";
    tmp(62000) := x"0800";
    tmp(62001) := x"0800";
    tmp(62002) := x"1000";
    tmp(62003) := x"1000";
    tmp(62004) := x"1000";
    tmp(62005) := x"1000";
    tmp(62006) := x"1000";
    tmp(62007) := x"1000";
    tmp(62008) := x"1000";
    tmp(62009) := x"1000";
    tmp(62010) := x"1000";
    tmp(62011) := x"1800";
    tmp(62012) := x"1800";
    tmp(62013) := x"1800";
    tmp(62014) := x"2000";
    tmp(62015) := x"2000";
    tmp(62016) := x"2800";
    tmp(62017) := x"2800";
    tmp(62018) := x"2800";
    tmp(62019) := x"2800";
    tmp(62020) := x"2000";
    tmp(62021) := x"2000";
    tmp(62022) := x"1800";
    tmp(62023) := x"1800";
    tmp(62024) := x"1000";
    tmp(62025) := x"1000";
    tmp(62026) := x"0800";
    tmp(62027) := x"1000";
    tmp(62028) := x"2000";
    tmp(62029) := x"3000";
    tmp(62030) := x"4000";
    tmp(62031) := x"4000";
    tmp(62032) := x"4000";
    tmp(62033) := x"4800";
    tmp(62034) := x"4800";
    tmp(62035) := x"4800";
    tmp(62036) := x"4000";
    tmp(62037) := x"4000";
    tmp(62038) := x"4000";
    tmp(62039) := x"4000";
    tmp(62040) := x"4800";
    tmp(62041) := x"4800";
    tmp(62042) := x"5000";
    tmp(62043) := x"5000";
    tmp(62044) := x"5000";
    tmp(62045) := x"5800";
    tmp(62046) := x"5800";
    tmp(62047) := x"5800";
    tmp(62048) := x"5800";
    tmp(62049) := x"5800";
    tmp(62050) := x"5800";
    tmp(62051) := x"6000";
    tmp(62052) := x"6800";
    tmp(62053) := x"6800";
    tmp(62054) := x"6800";
    tmp(62055) := x"6000";
    tmp(62056) := x"6000";
    tmp(62057) := x"6800";
    tmp(62058) := x"7800";
    tmp(62059) := x"9020";
    tmp(62060) := x"7000";
    tmp(62061) := x"6000";
    tmp(62062) := x"5800";
    tmp(62063) := x"6820";
    tmp(62064) := x"6820";
    tmp(62065) := x"6020";
    tmp(62066) := x"6020";
    tmp(62067) := x"6820";
    tmp(62068) := x"7020";
    tmp(62069) := x"6820";
    tmp(62070) := x"7020";
    tmp(62071) := x"9020";
    tmp(62072) := x"6820";
    tmp(62073) := x"6820";
    tmp(62074) := x"6820";
    tmp(62075) := x"8020";
    tmp(62076) := x"9020";
    tmp(62077) := x"9020";
    tmp(62078) := x"9820";
    tmp(62079) := x"a020";
    tmp(62080) := x"9020";
    tmp(62081) := x"9020";
    tmp(62082) := x"8020";
    tmp(62083) := x"9020";
    tmp(62084) := x"9820";
    tmp(62085) := x"9020";
    tmp(62086) := x"7800";
    tmp(62087) := x"7800";
    tmp(62088) := x"7800";
    tmp(62089) := x"8000";
    tmp(62090) := x"9000";
    tmp(62091) := x"9800";
    tmp(62092) := x"9800";
    tmp(62093) := x"8800";
    tmp(62094) := x"9800";
    tmp(62095) := x"a000";
    tmp(62096) := x"a820";
    tmp(62097) := x"b820";
    tmp(62098) := x"d020";
    tmp(62099) := x"8820";
    tmp(62100) := x"3841";
    tmp(62101) := x"1061";
    tmp(62102) := x"1081";
    tmp(62103) := x"1082";
    tmp(62104) := x"10a2";
    tmp(62105) := x"10a2";
    tmp(62106) := x"18a2";
    tmp(62107) := x"18a3";
    tmp(62108) := x"18c3";
    tmp(62109) := x"18c3";
    tmp(62110) := x"18c3";
    tmp(62111) := x"18c3";
    tmp(62112) := x"18c3";
    tmp(62113) := x"18c3";
    tmp(62114) := x"18c3";
    tmp(62115) := x"18e3";
    tmp(62116) := x"18e4";
    tmp(62117) := x"2104";
    tmp(62118) := x"2104";
    tmp(62119) := x"2104";
    tmp(62120) := x"2104";
    tmp(62121) := x"2104";
    tmp(62122) := x"2104";
    tmp(62123) := x"2125";
    tmp(62124) := x"2925";
    tmp(62125) := x"2925";
    tmp(62126) := x"2946";
    tmp(62127) := x"2946";
    tmp(62128) := x"2946";
    tmp(62129) := x"2966";
    tmp(62130) := x"2966";
    tmp(62131) := x"3166";
    tmp(62132) := x"3187";
    tmp(62133) := x"31a7";
    tmp(62134) := x"3187";
    tmp(62135) := x"31a8";
    tmp(62136) := x"39e8";
    tmp(62137) := x"39c8";
    tmp(62138) := x"39c8";
    tmp(62139) := x"39c8";
    tmp(62140) := x"41e9";
    tmp(62141) := x"420a";
    tmp(62142) := x"422a";
    tmp(62143) := x"422a";
    tmp(62144) := x"4a4b";
    tmp(62145) := x"4a4b";
    tmp(62146) := x"4a6b";
    tmp(62147) := x"4a4b";
    tmp(62148) := x"4a6b";
    tmp(62149) := x"4a8b";
    tmp(62150) := x"4a6b";
    tmp(62151) := x"4a6a";
    tmp(62152) := x"4a4a";
    tmp(62153) := x"4a4a";
    tmp(62154) := x"424a";
    tmp(62155) := x"4a4a";
    tmp(62156) := x"4a4a";
    tmp(62157) := x"424a";
    tmp(62158) := x"4249";
    tmp(62159) := x"3a28";
    tmp(62160) := x"0000";
    tmp(62161) := x"0800";
    tmp(62162) := x"0800";
    tmp(62163) := x"0800";
    tmp(62164) := x"0800";
    tmp(62165) := x"0800";
    tmp(62166) := x"1000";
    tmp(62167) := x"0800";
    tmp(62168) := x"1000";
    tmp(62169) := x"1000";
    tmp(62170) := x"1000";
    tmp(62171) := x"1000";
    tmp(62172) := x"1000";
    tmp(62173) := x"1000";
    tmp(62174) := x"1000";
    tmp(62175) := x"1000";
    tmp(62176) := x"1000";
    tmp(62177) := x"1000";
    tmp(62178) := x"1000";
    tmp(62179) := x"1000";
    tmp(62180) := x"1000";
    tmp(62181) := x"1000";
    tmp(62182) := x"1800";
    tmp(62183) := x"1800";
    tmp(62184) := x"1800";
    tmp(62185) := x"1000";
    tmp(62186) := x"1000";
    tmp(62187) := x"1000";
    tmp(62188) := x"1800";
    tmp(62189) := x"1800";
    tmp(62190) := x"1800";
    tmp(62191) := x"1800";
    tmp(62192) := x"1800";
    tmp(62193) := x"1800";
    tmp(62194) := x"2000";
    tmp(62195) := x"2000";
    tmp(62196) := x"1800";
    tmp(62197) := x"1800";
    tmp(62198) := x"1800";
    tmp(62199) := x"1800";
    tmp(62200) := x"1800";
    tmp(62201) := x"1800";
    tmp(62202) := x"2000";
    tmp(62203) := x"2000";
    tmp(62204) := x"2000";
    tmp(62205) := x"2800";
    tmp(62206) := x"2800";
    tmp(62207) := x"2800";
    tmp(62208) := x"2800";
    tmp(62209) := x"2000";
    tmp(62210) := x"2000";
    tmp(62211) := x"2000";
    tmp(62212) := x"2000";
    tmp(62213) := x"2000";
    tmp(62214) := x"2800";
    tmp(62215) := x"2800";
    tmp(62216) := x"2800";
    tmp(62217) := x"2800";
    tmp(62218) := x"3000";
    tmp(62219) := x"3000";
    tmp(62220) := x"3000";
    tmp(62221) := x"3000";
    tmp(62222) := x"3000";
    tmp(62223) := x"3000";
    tmp(62224) := x"3020";
    tmp(62225) := x"3020";
    tmp(62226) := x"2800";
    tmp(62227) := x"2000";
    tmp(62228) := x"1800";
    tmp(62229) := x"1800";
    tmp(62230) := x"1800";
    tmp(62231) := x"2000";
    tmp(62232) := x"2000";
    tmp(62233) := x"1800";
    tmp(62234) := x"1000";
    tmp(62235) := x"1000";
    tmp(62236) := x"1000";
    tmp(62237) := x"0820";
    tmp(62238) := x"0820";
    tmp(62239) := x"0800";
    tmp(62240) := x"0800";
    tmp(62241) := x"1000";
    tmp(62242) := x"1000";
    tmp(62243) := x"1000";
    tmp(62244) := x"1000";
    tmp(62245) := x"1000";
    tmp(62246) := x"0800";
    tmp(62247) := x"0800";
    tmp(62248) := x"0800";
    tmp(62249) := x"1000";
    tmp(62250) := x"1000";
    tmp(62251) := x"1800";
    tmp(62252) := x"2000";
    tmp(62253) := x"2800";
    tmp(62254) := x"3000";
    tmp(62255) := x"3000";
    tmp(62256) := x"3000";
    tmp(62257) := x"3000";
    tmp(62258) := x"2800";
    tmp(62259) := x"2000";
    tmp(62260) := x"2000";
    tmp(62261) := x"1800";
    tmp(62262) := x"1800";
    tmp(62263) := x"1800";
    tmp(62264) := x"1800";
    tmp(62265) := x"1000";
    tmp(62266) := x"1000";
    tmp(62267) := x"1800";
    tmp(62268) := x"2800";
    tmp(62269) := x"3000";
    tmp(62270) := x"3800";
    tmp(62271) := x"4000";
    tmp(62272) := x"4000";
    tmp(62273) := x"4000";
    tmp(62274) := x"4000";
    tmp(62275) := x"3800";
    tmp(62276) := x"3800";
    tmp(62277) := x"4000";
    tmp(62278) := x"4000";
    tmp(62279) := x"4000";
    tmp(62280) := x"4800";
    tmp(62281) := x"4800";
    tmp(62282) := x"4800";
    tmp(62283) := x"4800";
    tmp(62284) := x"5000";
    tmp(62285) := x"5800";
    tmp(62286) := x"5800";
    tmp(62287) := x"5000";
    tmp(62288) := x"5800";
    tmp(62289) := x"5800";
    tmp(62290) := x"5000";
    tmp(62291) := x"6000";
    tmp(62292) := x"6800";
    tmp(62293) := x"7000";
    tmp(62294) := x"7000";
    tmp(62295) := x"6000";
    tmp(62296) := x"6800";
    tmp(62297) := x"7000";
    tmp(62298) := x"8000";
    tmp(62299) := x"9020";
    tmp(62300) := x"6800";
    tmp(62301) := x"6000";
    tmp(62302) := x"5800";
    tmp(62303) := x"6820";
    tmp(62304) := x"6820";
    tmp(62305) := x"6020";
    tmp(62306) := x"6020";
    tmp(62307) := x"6820";
    tmp(62308) := x"7820";
    tmp(62309) := x"6820";
    tmp(62310) := x"7020";
    tmp(62311) := x"9840";
    tmp(62312) := x"7020";
    tmp(62313) := x"7020";
    tmp(62314) := x"7020";
    tmp(62315) := x"8820";
    tmp(62316) := x"9020";
    tmp(62317) := x"9820";
    tmp(62318) := x"a020";
    tmp(62319) := x"9820";
    tmp(62320) := x"8820";
    tmp(62321) := x"8020";
    tmp(62322) := x"8020";
    tmp(62323) := x"a840";
    tmp(62324) := x"9020";
    tmp(62325) := x"9020";
    tmp(62326) := x"8820";
    tmp(62327) := x"7800";
    tmp(62328) := x"7800";
    tmp(62329) := x"7800";
    tmp(62330) := x"8000";
    tmp(62331) := x"9000";
    tmp(62332) := x"9000";
    tmp(62333) := x"9000";
    tmp(62334) := x"9000";
    tmp(62335) := x"9800";
    tmp(62336) := x"a820";
    tmp(62337) := x"a800";
    tmp(62338) := x"c820";
    tmp(62339) := x"7020";
    tmp(62340) := x"2041";
    tmp(62341) := x"1061";
    tmp(62342) := x"1081";
    tmp(62343) := x"1082";
    tmp(62344) := x"10a2";
    tmp(62345) := x"10a2";
    tmp(62346) := x"10a2";
    tmp(62347) := x"18a2";
    tmp(62348) := x"18a3";
    tmp(62349) := x"18a2";
    tmp(62350) := x"18a3";
    tmp(62351) := x"18a3";
    tmp(62352) := x"18a3";
    tmp(62353) := x"18c3";
    tmp(62354) := x"18c3";
    tmp(62355) := x"18c3";
    tmp(62356) := x"18e3";
    tmp(62357) := x"18e3";
    tmp(62358) := x"20e4";
    tmp(62359) := x"2104";
    tmp(62360) := x"2104";
    tmp(62361) := x"2104";
    tmp(62362) := x"2104";
    tmp(62363) := x"2124";
    tmp(62364) := x"2125";
    tmp(62365) := x"2925";
    tmp(62366) := x"2925";
    tmp(62367) := x"2945";
    tmp(62368) := x"2125";
    tmp(62369) := x"2946";
    tmp(62370) := x"2946";
    tmp(62371) := x"2966";
    tmp(62372) := x"2966";
    tmp(62373) := x"3187";
    tmp(62374) := x"3187";
    tmp(62375) := x"31a7";
    tmp(62376) := x"39c7";
    tmp(62377) := x"39c7";
    tmp(62378) := x"39c8";
    tmp(62379) := x"39e8";
    tmp(62380) := x"41e9";
    tmp(62381) := x"41e9";
    tmp(62382) := x"4209";
    tmp(62383) := x"422a";
    tmp(62384) := x"4a4b";
    tmp(62385) := x"4a4a";
    tmp(62386) := x"4a6b";
    tmp(62387) := x"526b";
    tmp(62388) := x"52ac";
    tmp(62389) := x"52cd";
    tmp(62390) := x"52cd";
    tmp(62391) := x"52ac";
    tmp(62392) := x"528b";
    tmp(62393) := x"528b";
    tmp(62394) := x"528b";
    tmp(62395) := x"52ac";
    tmp(62396) := x"52ac";
    tmp(62397) := x"52ab";
    tmp(62398) := x"4a8b";
    tmp(62399) := x"426a";
    tmp(62400) := x"0000";
    tmp(62401) := x"0800";
    tmp(62402) := x"0800";
    tmp(62403) := x"0800";
    tmp(62404) := x"0800";
    tmp(62405) := x"0800";
    tmp(62406) := x"0800";
    tmp(62407) := x"0800";
    tmp(62408) := x"1000";
    tmp(62409) := x"1000";
    tmp(62410) := x"1000";
    tmp(62411) := x"1000";
    tmp(62412) := x"1000";
    tmp(62413) := x"1000";
    tmp(62414) := x"1000";
    tmp(62415) := x"1000";
    tmp(62416) := x"1000";
    tmp(62417) := x"1000";
    tmp(62418) := x"1000";
    tmp(62419) := x"1000";
    tmp(62420) := x"1000";
    tmp(62421) := x"1000";
    tmp(62422) := x"1000";
    tmp(62423) := x"1800";
    tmp(62424) := x"1000";
    tmp(62425) := x"1000";
    tmp(62426) := x"1000";
    tmp(62427) := x"1000";
    tmp(62428) := x"1000";
    tmp(62429) := x"1800";
    tmp(62430) := x"1800";
    tmp(62431) := x"1800";
    tmp(62432) := x"1800";
    tmp(62433) := x"2000";
    tmp(62434) := x"2000";
    tmp(62435) := x"2000";
    tmp(62436) := x"2000";
    tmp(62437) := x"2000";
    tmp(62438) := x"2000";
    tmp(62439) := x"1800";
    tmp(62440) := x"1800";
    tmp(62441) := x"1800";
    tmp(62442) := x"2000";
    tmp(62443) := x"2000";
    tmp(62444) := x"2000";
    tmp(62445) := x"2800";
    tmp(62446) := x"2800";
    tmp(62447) := x"2800";
    tmp(62448) := x"2800";
    tmp(62449) := x"2800";
    tmp(62450) := x"2000";
    tmp(62451) := x"2000";
    tmp(62452) := x"2000";
    tmp(62453) := x"2000";
    tmp(62454) := x"2800";
    tmp(62455) := x"2800";
    tmp(62456) := x"3000";
    tmp(62457) := x"3000";
    tmp(62458) := x"3000";
    tmp(62459) := x"3000";
    tmp(62460) := x"3800";
    tmp(62461) := x"3800";
    tmp(62462) := x"3800";
    tmp(62463) := x"3820";
    tmp(62464) := x"3000";
    tmp(62465) := x"2800";
    tmp(62466) := x"2800";
    tmp(62467) := x"2000";
    tmp(62468) := x"2000";
    tmp(62469) := x"2800";
    tmp(62470) := x"2800";
    tmp(62471) := x"2000";
    tmp(62472) := x"2000";
    tmp(62473) := x"1800";
    tmp(62474) := x"1800";
    tmp(62475) := x"1000";
    tmp(62476) := x"0800";
    tmp(62477) := x"0800";
    tmp(62478) := x"0800";
    tmp(62479) := x"0800";
    tmp(62480) := x"0800";
    tmp(62481) := x"0800";
    tmp(62482) := x"0800";
    tmp(62483) := x"0800";
    tmp(62484) := x"0800";
    tmp(62485) := x"0800";
    tmp(62486) := x"0800";
    tmp(62487) := x"0800";
    tmp(62488) := x"0800";
    tmp(62489) := x"1000";
    tmp(62490) := x"1000";
    tmp(62491) := x"1800";
    tmp(62492) := x"1800";
    tmp(62493) := x"2000";
    tmp(62494) := x"2800";
    tmp(62495) := x"2800";
    tmp(62496) := x"2800";
    tmp(62497) := x"2800";
    tmp(62498) := x"2800";
    tmp(62499) := x"2000";
    tmp(62500) := x"2000";
    tmp(62501) := x"1800";
    tmp(62502) := x"1800";
    tmp(62503) := x"1800";
    tmp(62504) := x"2000";
    tmp(62505) := x"2000";
    tmp(62506) := x"2000";
    tmp(62507) := x"2000";
    tmp(62508) := x"2800";
    tmp(62509) := x"3000";
    tmp(62510) := x"3000";
    tmp(62511) := x"3800";
    tmp(62512) := x"3800";
    tmp(62513) := x"3000";
    tmp(62514) := x"3000";
    tmp(62515) := x"3800";
    tmp(62516) := x"4000";
    tmp(62517) := x"4000";
    tmp(62518) := x"4000";
    tmp(62519) := x"4800";
    tmp(62520) := x"4800";
    tmp(62521) := x"4000";
    tmp(62522) := x"4800";
    tmp(62523) := x"5000";
    tmp(62524) := x"5000";
    tmp(62525) := x"5000";
    tmp(62526) := x"5000";
    tmp(62527) := x"5000";
    tmp(62528) := x"5800";
    tmp(62529) := x"5000";
    tmp(62530) := x"5000";
    tmp(62531) := x"6000";
    tmp(62532) := x"6800";
    tmp(62533) := x"7820";
    tmp(62534) := x"6800";
    tmp(62535) := x"6000";
    tmp(62536) := x"6800";
    tmp(62537) := x"8020";
    tmp(62538) := x"8020";
    tmp(62539) := x"8020";
    tmp(62540) := x"7000";
    tmp(62541) := x"7020";
    tmp(62542) := x"6020";
    tmp(62543) := x"6820";
    tmp(62544) := x"6820";
    tmp(62545) := x"5800";
    tmp(62546) := x"6020";
    tmp(62547) := x"6820";
    tmp(62548) := x"8840";
    tmp(62549) := x"7020";
    tmp(62550) := x"7820";
    tmp(62551) := x"9040";
    tmp(62552) := x"8820";
    tmp(62553) := x"7820";
    tmp(62554) := x"7820";
    tmp(62555) := x"8020";
    tmp(62556) := x"9020";
    tmp(62557) := x"9820";
    tmp(62558) := x"a020";
    tmp(62559) := x"a020";
    tmp(62560) := x"8820";
    tmp(62561) := x"7820";
    tmp(62562) := x"8820";
    tmp(62563) := x"b040";
    tmp(62564) := x"8820";
    tmp(62565) := x"8820";
    tmp(62566) := x"8820";
    tmp(62567) := x"7000";
    tmp(62568) := x"7800";
    tmp(62569) := x"7000";
    tmp(62570) := x"7800";
    tmp(62571) := x"9000";
    tmp(62572) := x"9000";
    tmp(62573) := x"8800";
    tmp(62574) := x"9000";
    tmp(62575) := x"9000";
    tmp(62576) := x"a000";
    tmp(62577) := x"9800";
    tmp(62578) := x"b820";
    tmp(62579) := x"5040";
    tmp(62580) := x"1041";
    tmp(62581) := x"1061";
    tmp(62582) := x"1081";
    tmp(62583) := x"1081";
    tmp(62584) := x"1082";
    tmp(62585) := x"10a2";
    tmp(62586) := x"10a2";
    tmp(62587) := x"10a2";
    tmp(62588) := x"10a2";
    tmp(62589) := x"10a2";
    tmp(62590) := x"10a2";
    tmp(62591) := x"10a2";
    tmp(62592) := x"10a2";
    tmp(62593) := x"10a2";
    tmp(62594) := x"18c3";
    tmp(62595) := x"18a3";
    tmp(62596) := x"18c3";
    tmp(62597) := x"18c3";
    tmp(62598) := x"18e3";
    tmp(62599) := x"18e3";
    tmp(62600) := x"20e4";
    tmp(62601) := x"2104";
    tmp(62602) := x"2104";
    tmp(62603) := x"2104";
    tmp(62604) := x"2104";
    tmp(62605) := x"2104";
    tmp(62606) := x"2104";
    tmp(62607) := x"2104";
    tmp(62608) := x"2125";
    tmp(62609) := x"2125";
    tmp(62610) := x"2945";
    tmp(62611) := x"2945";
    tmp(62612) := x"2966";
    tmp(62613) := x"3166";
    tmp(62614) := x"31a7";
    tmp(62615) := x"31a7";
    tmp(62616) := x"31a7";
    tmp(62617) := x"39a7";
    tmp(62618) := x"39c8";
    tmp(62619) := x"39e8";
    tmp(62620) := x"41e9";
    tmp(62621) := x"420a";
    tmp(62622) := x"422a";
    tmp(62623) := x"4a4b";
    tmp(62624) := x"4a4b";
    tmp(62625) := x"526b";
    tmp(62626) := x"528c";
    tmp(62627) := x"5aad";
    tmp(62628) := x"5aee";
    tmp(62629) := x"632f";
    tmp(62630) := x"632f";
    tmp(62631) := x"5b0e";
    tmp(62632) := x"5acd";
    tmp(62633) := x"5acd";
    tmp(62634) := x"5acd";
    tmp(62635) := x"5acd";
    tmp(62636) := x"5aed";
    tmp(62637) := x"5acd";
    tmp(62638) := x"52ab";
    tmp(62639) := x"4a8b";
    tmp(62640) := x"0000";
    tmp(62641) := x"0800";
    tmp(62642) := x"0800";
    tmp(62643) := x"0800";
    tmp(62644) := x"0800";
    tmp(62645) := x"0800";
    tmp(62646) := x"0800";
    tmp(62647) := x"1000";
    tmp(62648) := x"1000";
    tmp(62649) := x"1000";
    tmp(62650) := x"1000";
    tmp(62651) := x"1000";
    tmp(62652) := x"1000";
    tmp(62653) := x"1000";
    tmp(62654) := x"1000";
    tmp(62655) := x"1000";
    tmp(62656) := x"1000";
    tmp(62657) := x"1000";
    tmp(62658) := x"1000";
    tmp(62659) := x"1000";
    tmp(62660) := x"1000";
    tmp(62661) := x"1000";
    tmp(62662) := x"1800";
    tmp(62663) := x"1800";
    tmp(62664) := x"1000";
    tmp(62665) := x"1000";
    tmp(62666) := x"1000";
    tmp(62667) := x"1000";
    tmp(62668) := x"1000";
    tmp(62669) := x"1800";
    tmp(62670) := x"1800";
    tmp(62671) := x"1800";
    tmp(62672) := x"1800";
    tmp(62673) := x"2000";
    tmp(62674) := x"2000";
    tmp(62675) := x"2000";
    tmp(62676) := x"2000";
    tmp(62677) := x"2000";
    tmp(62678) := x"2000";
    tmp(62679) := x"1800";
    tmp(62680) := x"1800";
    tmp(62681) := x"2000";
    tmp(62682) := x"2000";
    tmp(62683) := x"2000";
    tmp(62684) := x"2000";
    tmp(62685) := x"2000";
    tmp(62686) := x"2800";
    tmp(62687) := x"2800";
    tmp(62688) := x"2800";
    tmp(62689) := x"2000";
    tmp(62690) := x"2000";
    tmp(62691) := x"2000";
    tmp(62692) := x"2000";
    tmp(62693) := x"2800";
    tmp(62694) := x"2800";
    tmp(62695) := x"2800";
    tmp(62696) := x"2800";
    tmp(62697) := x"3000";
    tmp(62698) := x"3000";
    tmp(62699) := x"3800";
    tmp(62700) := x"3800";
    tmp(62701) := x"3800";
    tmp(62702) := x"3800";
    tmp(62703) := x"3000";
    tmp(62704) := x"3000";
    tmp(62705) := x"2800";
    tmp(62706) := x"2800";
    tmp(62707) := x"2800";
    tmp(62708) := x"2800";
    tmp(62709) := x"2800";
    tmp(62710) := x"2800";
    tmp(62711) := x"2000";
    tmp(62712) := x"2000";
    tmp(62713) := x"1800";
    tmp(62714) := x"1000";
    tmp(62715) := x"1000";
    tmp(62716) := x"0800";
    tmp(62717) := x"0800";
    tmp(62718) := x"0800";
    tmp(62719) := x"0800";
    tmp(62720) := x"1000";
    tmp(62721) := x"0800";
    tmp(62722) := x"0800";
    tmp(62723) := x"0800";
    tmp(62724) := x"0820";
    tmp(62725) := x"0800";
    tmp(62726) := x"0800";
    tmp(62727) := x"0800";
    tmp(62728) := x"0800";
    tmp(62729) := x"1000";
    tmp(62730) := x"1000";
    tmp(62731) := x"1000";
    tmp(62732) := x"1800";
    tmp(62733) := x"1800";
    tmp(62734) := x"1800";
    tmp(62735) := x"1800";
    tmp(62736) := x"1800";
    tmp(62737) := x"1800";
    tmp(62738) := x"1800";
    tmp(62739) := x"1800";
    tmp(62740) := x"1800";
    tmp(62741) := x"1800";
    tmp(62742) := x"1800";
    tmp(62743) := x"1800";
    tmp(62744) := x"1800";
    tmp(62745) := x"1000";
    tmp(62746) := x"1000";
    tmp(62747) := x"2000";
    tmp(62748) := x"2800";
    tmp(62749) := x"2800";
    tmp(62750) := x"2800";
    tmp(62751) := x"2800";
    tmp(62752) := x"2800";
    tmp(62753) := x"2800";
    tmp(62754) := x"3000";
    tmp(62755) := x"3800";
    tmp(62756) := x"3800";
    tmp(62757) := x"3800";
    tmp(62758) := x"4800";
    tmp(62759) := x"4800";
    tmp(62760) := x"4000";
    tmp(62761) := x"4800";
    tmp(62762) := x"5000";
    tmp(62763) := x"5000";
    tmp(62764) := x"5000";
    tmp(62765) := x"5000";
    tmp(62766) := x"5000";
    tmp(62767) := x"5000";
    tmp(62768) := x"5800";
    tmp(62769) := x"5000";
    tmp(62770) := x"5000";
    tmp(62771) := x"6800";
    tmp(62772) := x"6800";
    tmp(62773) := x"7000";
    tmp(62774) := x"7000";
    tmp(62775) := x"6800";
    tmp(62776) := x"6800";
    tmp(62777) := x"7000";
    tmp(62778) := x"7800";
    tmp(62779) := x"8020";
    tmp(62780) := x"7820";
    tmp(62781) := x"6820";
    tmp(62782) := x"5800";
    tmp(62783) := x"6020";
    tmp(62784) := x"6020";
    tmp(62785) := x"6020";
    tmp(62786) := x"5800";
    tmp(62787) := x"7820";
    tmp(62788) := x"9040";
    tmp(62789) := x"7820";
    tmp(62790) := x"8020";
    tmp(62791) := x"9020";
    tmp(62792) := x"8820";
    tmp(62793) := x"7820";
    tmp(62794) := x"7020";
    tmp(62795) := x"8020";
    tmp(62796) := x"9820";
    tmp(62797) := x"9820";
    tmp(62798) := x"a820";
    tmp(62799) := x"9020";
    tmp(62800) := x"8020";
    tmp(62801) := x"7820";
    tmp(62802) := x"8820";
    tmp(62803) := x"a840";
    tmp(62804) := x"8820";
    tmp(62805) := x"9020";
    tmp(62806) := x"8820";
    tmp(62807) := x"7000";
    tmp(62808) := x"7000";
    tmp(62809) := x"7000";
    tmp(62810) := x"7800";
    tmp(62811) := x"8800";
    tmp(62812) := x"9020";
    tmp(62813) := x"8800";
    tmp(62814) := x"9820";
    tmp(62815) := x"9000";
    tmp(62816) := x"9000";
    tmp(62817) := x"9800";
    tmp(62818) := x"9820";
    tmp(62819) := x"3041";
    tmp(62820) := x"1061";
    tmp(62821) := x"1061";
    tmp(62822) := x"1081";
    tmp(62823) := x"1081";
    tmp(62824) := x"1082";
    tmp(62825) := x"1082";
    tmp(62826) := x"1082";
    tmp(62827) := x"1082";
    tmp(62828) := x"1082";
    tmp(62829) := x"1082";
    tmp(62830) := x"1082";
    tmp(62831) := x"1082";
    tmp(62832) := x"1082";
    tmp(62833) := x"10a2";
    tmp(62834) := x"10a2";
    tmp(62835) := x"10a2";
    tmp(62836) := x"18a2";
    tmp(62837) := x"18c3";
    tmp(62838) := x"18e3";
    tmp(62839) := x"18e3";
    tmp(62840) := x"18e3";
    tmp(62841) := x"20e3";
    tmp(62842) := x"20e3";
    tmp(62843) := x"20e3";
    tmp(62844) := x"20e3";
    tmp(62845) := x"2103";
    tmp(62846) := x"2104";
    tmp(62847) := x"2104";
    tmp(62848) := x"2104";
    tmp(62849) := x"2105";
    tmp(62850) := x"2125";
    tmp(62851) := x"2945";
    tmp(62852) := x"2966";
    tmp(62853) := x"3186";
    tmp(62854) := x"3186";
    tmp(62855) := x"39a7";
    tmp(62856) := x"39a7";
    tmp(62857) := x"39c8";
    tmp(62858) := x"41e8";
    tmp(62859) := x"4209";
    tmp(62860) := x"4a09";
    tmp(62861) := x"4a2a";
    tmp(62862) := x"4a4b";
    tmp(62863) := x"528c";
    tmp(62864) := x"5acd";
    tmp(62865) := x"62ce";
    tmp(62866) := x"62ee";
    tmp(62867) := x"630f";
    tmp(62868) := x"6b50";
    tmp(62869) := x"7371";
    tmp(62870) := x"7371";
    tmp(62871) := x"6b50";
    tmp(62872) := x"632f";
    tmp(62873) := x"632f";
    tmp(62874) := x"630f";
    tmp(62875) := x"630f";
    tmp(62876) := x"632e";
    tmp(62877) := x"5b0e";
    tmp(62878) := x"52ed";
    tmp(62879) := x"52cc";
    tmp(62880) := x"0000";
    tmp(62881) := x"0800";
    tmp(62882) := x"0800";
    tmp(62883) := x"0800";
    tmp(62884) := x"0800";
    tmp(62885) := x"0800";
    tmp(62886) := x"0800";
    tmp(62887) := x"1000";
    tmp(62888) := x"1000";
    tmp(62889) := x"1000";
    tmp(62890) := x"1000";
    tmp(62891) := x"1000";
    tmp(62892) := x"1000";
    tmp(62893) := x"1000";
    tmp(62894) := x"1000";
    tmp(62895) := x"1000";
    tmp(62896) := x"1000";
    tmp(62897) := x"1000";
    tmp(62898) := x"1000";
    tmp(62899) := x"1000";
    tmp(62900) := x"1000";
    tmp(62901) := x"1000";
    tmp(62902) := x"1000";
    tmp(62903) := x"1800";
    tmp(62904) := x"1800";
    tmp(62905) := x"1000";
    tmp(62906) := x"1000";
    tmp(62907) := x"1000";
    tmp(62908) := x"1000";
    tmp(62909) := x"1800";
    tmp(62910) := x"1800";
    tmp(62911) := x"1800";
    tmp(62912) := x"1800";
    tmp(62913) := x"1800";
    tmp(62914) := x"2000";
    tmp(62915) := x"2000";
    tmp(62916) := x"2000";
    tmp(62917) := x"2000";
    tmp(62918) := x"2000";
    tmp(62919) := x"1800";
    tmp(62920) := x"2000";
    tmp(62921) := x"2000";
    tmp(62922) := x"2000";
    tmp(62923) := x"2000";
    tmp(62924) := x"2800";
    tmp(62925) := x"2800";
    tmp(62926) := x"2800";
    tmp(62927) := x"2800";
    tmp(62928) := x"2800";
    tmp(62929) := x"2000";
    tmp(62930) := x"2000";
    tmp(62931) := x"2000";
    tmp(62932) := x"2000";
    tmp(62933) := x"2800";
    tmp(62934) := x"2800";
    tmp(62935) := x"2800";
    tmp(62936) := x"2800";
    tmp(62937) := x"2800";
    tmp(62938) := x"3000";
    tmp(62939) := x"3000";
    tmp(62940) := x"3000";
    tmp(62941) := x"3000";
    tmp(62942) := x"3000";
    tmp(62943) := x"3000";
    tmp(62944) := x"3000";
    tmp(62945) := x"3000";
    tmp(62946) := x"3000";
    tmp(62947) := x"2800";
    tmp(62948) := x"2800";
    tmp(62949) := x"2800";
    tmp(62950) := x"2000";
    tmp(62951) := x"2000";
    tmp(62952) := x"2000";
    tmp(62953) := x"1800";
    tmp(62954) := x"1000";
    tmp(62955) := x"0800";
    tmp(62956) := x"0800";
    tmp(62957) := x"0800";
    tmp(62958) := x"0800";
    tmp(62959) := x"1000";
    tmp(62960) := x"1000";
    tmp(62961) := x"1000";
    tmp(62962) := x"1020";
    tmp(62963) := x"0820";
    tmp(62964) := x"0820";
    tmp(62965) := x"0820";
    tmp(62966) := x"0820";
    tmp(62967) := x"0800";
    tmp(62968) := x"1000";
    tmp(62969) := x"1000";
    tmp(62970) := x"1000";
    tmp(62971) := x"1000";
    tmp(62972) := x"1000";
    tmp(62973) := x"1800";
    tmp(62974) := x"1800";
    tmp(62975) := x"1800";
    tmp(62976) := x"1800";
    tmp(62977) := x"1800";
    tmp(62978) := x"1800";
    tmp(62979) := x"1800";
    tmp(62980) := x"1800";
    tmp(62981) := x"1000";
    tmp(62982) := x"1000";
    tmp(62983) := x"1000";
    tmp(62984) := x"1000";
    tmp(62985) := x"1000";
    tmp(62986) := x"1000";
    tmp(62987) := x"1800";
    tmp(62988) := x"2000";
    tmp(62989) := x"2000";
    tmp(62990) := x"1800";
    tmp(62991) := x"1800";
    tmp(62992) := x"2000";
    tmp(62993) := x"3000";
    tmp(62994) := x"3800";
    tmp(62995) := x"3800";
    tmp(62996) := x"3800";
    tmp(62997) := x"4000";
    tmp(62998) := x"4800";
    tmp(62999) := x"4000";
    tmp(63000) := x"4800";
    tmp(63001) := x"4800";
    tmp(63002) := x"5000";
    tmp(63003) := x"5000";
    tmp(63004) := x"5800";
    tmp(63005) := x"5800";
    tmp(63006) := x"5800";
    tmp(63007) := x"5800";
    tmp(63008) := x"5800";
    tmp(63009) := x"5000";
    tmp(63010) := x"5800";
    tmp(63011) := x"6000";
    tmp(63012) := x"6000";
    tmp(63013) := x"6800";
    tmp(63014) := x"6800";
    tmp(63015) := x"7000";
    tmp(63016) := x"6800";
    tmp(63017) := x"6800";
    tmp(63018) := x"7800";
    tmp(63019) := x"8020";
    tmp(63020) := x"6800";
    tmp(63021) := x"6000";
    tmp(63022) := x"5000";
    tmp(63023) := x"6020";
    tmp(63024) := x"5800";
    tmp(63025) := x"5800";
    tmp(63026) := x"6000";
    tmp(63027) := x"7020";
    tmp(63028) := x"8820";
    tmp(63029) := x"7820";
    tmp(63030) := x"7820";
    tmp(63031) := x"9020";
    tmp(63032) := x"8020";
    tmp(63033) := x"7820";
    tmp(63034) := x"8020";
    tmp(63035) := x"8820";
    tmp(63036) := x"9020";
    tmp(63037) := x"8820";
    tmp(63038) := x"9820";
    tmp(63039) := x"8820";
    tmp(63040) := x"8020";
    tmp(63041) := x"8020";
    tmp(63042) := x"8020";
    tmp(63043) := x"b040";
    tmp(63044) := x"9020";
    tmp(63045) := x"9020";
    tmp(63046) := x"9020";
    tmp(63047) := x"7800";
    tmp(63048) := x"6800";
    tmp(63049) := x"7000";
    tmp(63050) := x"8800";
    tmp(63051) := x"8820";
    tmp(63052) := x"8820";
    tmp(63053) := x"8820";
    tmp(63054) := x"9020";
    tmp(63055) := x"8800";
    tmp(63056) := x"8800";
    tmp(63057) := x"9000";
    tmp(63058) := x"7820";
    tmp(63059) := x"2041";
    tmp(63060) := x"1061";
    tmp(63061) := x"1061";
    tmp(63062) := x"1061";
    tmp(63063) := x"1061";
    tmp(63064) := x"1081";
    tmp(63065) := x"1081";
    tmp(63066) := x"1082";
    tmp(63067) := x"1082";
    tmp(63068) := x"1082";
    tmp(63069) := x"1082";
    tmp(63070) := x"1082";
    tmp(63071) := x"1081";
    tmp(63072) := x"1082";
    tmp(63073) := x"1082";
    tmp(63074) := x"1082";
    tmp(63075) := x"10a2";
    tmp(63076) := x"10a2";
    tmp(63077) := x"10a2";
    tmp(63078) := x"18c3";
    tmp(63079) := x"18c3";
    tmp(63080) := x"18e3";
    tmp(63081) := x"20e3";
    tmp(63082) := x"20e3";
    tmp(63083) := x"18e3";
    tmp(63084) := x"18e3";
    tmp(63085) := x"20e3";
    tmp(63086) := x"20e4";
    tmp(63087) := x"2104";
    tmp(63088) := x"2104";
    tmp(63089) := x"2104";
    tmp(63090) := x"2925";
    tmp(63091) := x"2966";
    tmp(63092) := x"3186";
    tmp(63093) := x"31a7";
    tmp(63094) := x"39a7";
    tmp(63095) := x"39c7";
    tmp(63096) := x"41e8";
    tmp(63097) := x"4209";
    tmp(63098) := x"4a2a";
    tmp(63099) := x"4a2a";
    tmp(63100) := x"524b";
    tmp(63101) := x"528c";
    tmp(63102) := x"5aee";
    tmp(63103) := x"5acd";
    tmp(63104) := x"630f";
    tmp(63105) := x"6310";
    tmp(63106) := x"7371";
    tmp(63107) := x"7372";
    tmp(63108) := x"73b2";
    tmp(63109) := x"7bd3";
    tmp(63110) := x"73b2";
    tmp(63111) := x"7392";
    tmp(63112) := x"7391";
    tmp(63113) := x"6b71";
    tmp(63114) := x"6b50";
    tmp(63115) := x"6b50";
    tmp(63116) := x"6b6f";
    tmp(63117) := x"634f";
    tmp(63118) := x"5b2e";
    tmp(63119) := x"5aed";
    tmp(63120) := x"0000";
    tmp(63121) := x"0800";
    tmp(63122) := x"0800";
    tmp(63123) := x"0800";
    tmp(63124) := x"0800";
    tmp(63125) := x"0800";
    tmp(63126) := x"0800";
    tmp(63127) := x"1000";
    tmp(63128) := x"1000";
    tmp(63129) := x"1000";
    tmp(63130) := x"1000";
    tmp(63131) := x"1000";
    tmp(63132) := x"1000";
    tmp(63133) := x"1000";
    tmp(63134) := x"1000";
    tmp(63135) := x"1000";
    tmp(63136) := x"1000";
    tmp(63137) := x"1000";
    tmp(63138) := x"1000";
    tmp(63139) := x"1000";
    tmp(63140) := x"1000";
    tmp(63141) := x"1000";
    tmp(63142) := x"1000";
    tmp(63143) := x"1000";
    tmp(63144) := x"1000";
    tmp(63145) := x"1000";
    tmp(63146) := x"1000";
    tmp(63147) := x"1000";
    tmp(63148) := x"1000";
    tmp(63149) := x"1000";
    tmp(63150) := x"1000";
    tmp(63151) := x"1800";
    tmp(63152) := x"1800";
    tmp(63153) := x"1800";
    tmp(63154) := x"1800";
    tmp(63155) := x"1800";
    tmp(63156) := x"1800";
    tmp(63157) := x"1800";
    tmp(63158) := x"1800";
    tmp(63159) := x"2000";
    tmp(63160) := x"2000";
    tmp(63161) := x"2000";
    tmp(63162) := x"2000";
    tmp(63163) := x"2000";
    tmp(63164) := x"2800";
    tmp(63165) := x"2800";
    tmp(63166) := x"2800";
    tmp(63167) := x"2800";
    tmp(63168) := x"2800";
    tmp(63169) := x"2800";
    tmp(63170) := x"2000";
    tmp(63171) := x"2000";
    tmp(63172) := x"2000";
    tmp(63173) := x"2000";
    tmp(63174) := x"2000";
    tmp(63175) := x"2800";
    tmp(63176) := x"2800";
    tmp(63177) := x"2800";
    tmp(63178) := x"2800";
    tmp(63179) := x"3000";
    tmp(63180) := x"3000";
    tmp(63181) := x"3000";
    tmp(63182) := x"3000";
    tmp(63183) := x"3000";
    tmp(63184) := x"3000";
    tmp(63185) := x"3000";
    tmp(63186) := x"2800";
    tmp(63187) := x"2800";
    tmp(63188) := x"2000";
    tmp(63189) := x"2000";
    tmp(63190) := x"2000";
    tmp(63191) := x"2000";
    tmp(63192) := x"1800";
    tmp(63193) := x"1000";
    tmp(63194) := x"0800";
    tmp(63195) := x"0800";
    tmp(63196) := x"0800";
    tmp(63197) := x"0800";
    tmp(63198) := x"1000";
    tmp(63199) := x"1000";
    tmp(63200) := x"1000";
    tmp(63201) := x"1000";
    tmp(63202) := x"1020";
    tmp(63203) := x"0820";
    tmp(63204) := x"0820";
    tmp(63205) := x"0820";
    tmp(63206) := x"1020";
    tmp(63207) := x"1020";
    tmp(63208) := x"0800";
    tmp(63209) := x"1000";
    tmp(63210) := x"1000";
    tmp(63211) := x"1000";
    tmp(63212) := x"1000";
    tmp(63213) := x"1000";
    tmp(63214) := x"1000";
    tmp(63215) := x"1000";
    tmp(63216) := x"0800";
    tmp(63217) := x"0800";
    tmp(63218) := x"0800";
    tmp(63219) := x"1000";
    tmp(63220) := x"1000";
    tmp(63221) := x"1800";
    tmp(63222) := x"1800";
    tmp(63223) := x"1800";
    tmp(63224) := x"1800";
    tmp(63225) := x"1800";
    tmp(63226) := x"1800";
    tmp(63227) := x"2000";
    tmp(63228) := x"2800";
    tmp(63229) := x"2000";
    tmp(63230) := x"1000";
    tmp(63231) := x"1800";
    tmp(63232) := x"2800";
    tmp(63233) := x"3000";
    tmp(63234) := x"3000";
    tmp(63235) := x"3800";
    tmp(63236) := x"3800";
    tmp(63237) := x"4000";
    tmp(63238) := x"3800";
    tmp(63239) := x"3800";
    tmp(63240) := x"4800";
    tmp(63241) := x"5000";
    tmp(63242) := x"5000";
    tmp(63243) := x"5000";
    tmp(63244) := x"5000";
    tmp(63245) := x"5800";
    tmp(63246) := x"6000";
    tmp(63247) := x"6000";
    tmp(63248) := x"5800";
    tmp(63249) := x"5800";
    tmp(63250) := x"6000";
    tmp(63251) := x"6000";
    tmp(63252) := x"6000";
    tmp(63253) := x"5800";
    tmp(63254) := x"6800";
    tmp(63255) := x"6800";
    tmp(63256) := x"6800";
    tmp(63257) := x"6800";
    tmp(63258) := x"7800";
    tmp(63259) := x"7800";
    tmp(63260) := x"6800";
    tmp(63261) := x"5800";
    tmp(63262) := x"5800";
    tmp(63263) := x"6820";
    tmp(63264) := x"5800";
    tmp(63265) := x"5000";
    tmp(63266) := x"6000";
    tmp(63267) := x"7020";
    tmp(63268) := x"8820";
    tmp(63269) := x"7820";
    tmp(63270) := x"7820";
    tmp(63271) := x"a020";
    tmp(63272) := x"8020";
    tmp(63273) := x"8020";
    tmp(63274) := x"7820";
    tmp(63275) := x"7820";
    tmp(63276) := x"8820";
    tmp(63277) := x"8820";
    tmp(63278) := x"9820";
    tmp(63279) := x"8820";
    tmp(63280) := x"8020";
    tmp(63281) := x"8820";
    tmp(63282) := x"7820";
    tmp(63283) := x"9820";
    tmp(63284) := x"8020";
    tmp(63285) := x"d061";
    tmp(63286) := x"8020";
    tmp(63287) := x"7800";
    tmp(63288) := x"7000";
    tmp(63289) := x"8020";
    tmp(63290) := x"9020";
    tmp(63291) := x"9020";
    tmp(63292) := x"8820";
    tmp(63293) := x"7800";
    tmp(63294) := x"9020";
    tmp(63295) := x"9000";
    tmp(63296) := x"8000";
    tmp(63297) := x"8800";
    tmp(63298) := x"5820";
    tmp(63299) := x"1041";
    tmp(63300) := x"1061";
    tmp(63301) := x"0861";
    tmp(63302) := x"1061";
    tmp(63303) := x"1061";
    tmp(63304) := x"1061";
    tmp(63305) := x"1061";
    tmp(63306) := x"1061";
    tmp(63307) := x"0861";
    tmp(63308) := x"1061";
    tmp(63309) := x"1061";
    tmp(63310) := x"1061";
    tmp(63311) := x"1061";
    tmp(63312) := x"1061";
    tmp(63313) := x"1081";
    tmp(63314) := x"1082";
    tmp(63315) := x"1082";
    tmp(63316) := x"10a2";
    tmp(63317) := x"18a2";
    tmp(63318) := x"18c3";
    tmp(63319) := x"18c3";
    tmp(63320) := x"20e3";
    tmp(63321) := x"2103";
    tmp(63322) := x"2104";
    tmp(63323) := x"20e3";
    tmp(63324) := x"20e3";
    tmp(63325) := x"20e4";
    tmp(63326) := x"2104";
    tmp(63327) := x"2124";
    tmp(63328) := x"2125";
    tmp(63329) := x"2945";
    tmp(63330) := x"2966";
    tmp(63331) := x"3186";
    tmp(63332) := x"39a7";
    tmp(63333) := x"39e8";
    tmp(63334) := x"41e8";
    tmp(63335) := x"41e9";
    tmp(63336) := x"422a";
    tmp(63337) := x"4a4a";
    tmp(63338) := x"524b";
    tmp(63339) := x"526c";
    tmp(63340) := x"5aad";
    tmp(63341) := x"630e";
    tmp(63342) := x"632e";
    tmp(63343) := x"6b2f";
    tmp(63344) := x"7371";
    tmp(63345) := x"7392";
    tmp(63346) := x"7bb3";
    tmp(63347) := x"8415";
    tmp(63348) := x"8c35";
    tmp(63349) := x"8c35";
    tmp(63350) := x"8435";
    tmp(63351) := x"83f4";
    tmp(63352) := x"7bf4";
    tmp(63353) := x"73b2";
    tmp(63354) := x"73b2";
    tmp(63355) := x"7371";
    tmp(63356) := x"7391";
    tmp(63357) := x"6b4f";
    tmp(63358) := x"634f";
    tmp(63359) := x"632f";
    tmp(63360) := x"0000";
    tmp(63361) := x"0800";
    tmp(63362) := x"0800";
    tmp(63363) := x"0800";
    tmp(63364) := x"0800";
    tmp(63365) := x"0800";
    tmp(63366) := x"1000";
    tmp(63367) := x"1000";
    tmp(63368) := x"1000";
    tmp(63369) := x"1000";
    tmp(63370) := x"1000";
    tmp(63371) := x"1000";
    tmp(63372) := x"1000";
    tmp(63373) := x"1000";
    tmp(63374) := x"1000";
    tmp(63375) := x"1000";
    tmp(63376) := x"1000";
    tmp(63377) := x"1000";
    tmp(63378) := x"1000";
    tmp(63379) := x"1000";
    tmp(63380) := x"1000";
    tmp(63381) := x"1000";
    tmp(63382) := x"1000";
    tmp(63383) := x"1000";
    tmp(63384) := x"1000";
    tmp(63385) := x"1000";
    tmp(63386) := x"1000";
    tmp(63387) := x"1000";
    tmp(63388) := x"1000";
    tmp(63389) := x"1000";
    tmp(63390) := x"1800";
    tmp(63391) := x"1800";
    tmp(63392) := x"1800";
    tmp(63393) := x"1800";
    tmp(63394) := x"1800";
    tmp(63395) := x"1800";
    tmp(63396) := x"1800";
    tmp(63397) := x"1800";
    tmp(63398) := x"1800";
    tmp(63399) := x"2000";
    tmp(63400) := x"2000";
    tmp(63401) := x"2000";
    tmp(63402) := x"2000";
    tmp(63403) := x"2000";
    tmp(63404) := x"2800";
    tmp(63405) := x"2800";
    tmp(63406) := x"2800";
    tmp(63407) := x"2800";
    tmp(63408) := x"2800";
    tmp(63409) := x"2800";
    tmp(63410) := x"2800";
    tmp(63411) := x"2000";
    tmp(63412) := x"2000";
    tmp(63413) := x"2000";
    tmp(63414) := x"2800";
    tmp(63415) := x"2800";
    tmp(63416) := x"2000";
    tmp(63417) := x"2800";
    tmp(63418) := x"2800";
    tmp(63419) := x"2800";
    tmp(63420) := x"2800";
    tmp(63421) := x"2800";
    tmp(63422) := x"3000";
    tmp(63423) := x"3000";
    tmp(63424) := x"2800";
    tmp(63425) := x"2800";
    tmp(63426) := x"2800";
    tmp(63427) := x"2800";
    tmp(63428) := x"2800";
    tmp(63429) := x"2000";
    tmp(63430) := x"2000";
    tmp(63431) := x"2000";
    tmp(63432) := x"1800";
    tmp(63433) := x"1000";
    tmp(63434) := x"1020";
    tmp(63435) := x"1020";
    tmp(63436) := x"0800";
    tmp(63437) := x"1000";
    tmp(63438) := x"1000";
    tmp(63439) := x"1000";
    tmp(63440) := x"1000";
    tmp(63441) := x"1000";
    tmp(63442) := x"1000";
    tmp(63443) := x"1020";
    tmp(63444) := x"1020";
    tmp(63445) := x"1020";
    tmp(63446) := x"0820";
    tmp(63447) := x"0820";
    tmp(63448) := x"0800";
    tmp(63449) := x"0800";
    tmp(63450) := x"0800";
    tmp(63451) := x"0800";
    tmp(63452) := x"0800";
    tmp(63453) := x"0800";
    tmp(63454) := x"0800";
    tmp(63455) := x"0800";
    tmp(63456) := x"1000";
    tmp(63457) := x"0800";
    tmp(63458) := x"0800";
    tmp(63459) := x"1000";
    tmp(63460) := x"1000";
    tmp(63461) := x"1000";
    tmp(63462) := x"0800";
    tmp(63463) := x"1000";
    tmp(63464) := x"1800";
    tmp(63465) := x"2000";
    tmp(63466) := x"2800";
    tmp(63467) := x"2000";
    tmp(63468) := x"1800";
    tmp(63469) := x"1000";
    tmp(63470) := x"1000";
    tmp(63471) := x"1800";
    tmp(63472) := x"2800";
    tmp(63473) := x"2800";
    tmp(63474) := x"2800";
    tmp(63475) := x"2800";
    tmp(63476) := x"2800";
    tmp(63477) := x"3800";
    tmp(63478) := x"3800";
    tmp(63479) := x"4000";
    tmp(63480) := x"4800";
    tmp(63481) := x"4800";
    tmp(63482) := x"5000";
    tmp(63483) := x"5800";
    tmp(63484) := x"5800";
    tmp(63485) := x"6000";
    tmp(63486) := x"6000";
    tmp(63487) := x"5800";
    tmp(63488) := x"5000";
    tmp(63489) := x"6000";
    tmp(63490) := x"6000";
    tmp(63491) := x"5800";
    tmp(63492) := x"6000";
    tmp(63493) := x"5800";
    tmp(63494) := x"6000";
    tmp(63495) := x"6000";
    tmp(63496) := x"6000";
    tmp(63497) := x"6800";
    tmp(63498) := x"8000";
    tmp(63499) := x"7000";
    tmp(63500) := x"6800";
    tmp(63501) := x"6000";
    tmp(63502) := x"6000";
    tmp(63503) := x"6820";
    tmp(63504) := x"6000";
    tmp(63505) := x"5800";
    tmp(63506) := x"6000";
    tmp(63507) := x"7020";
    tmp(63508) := x"8820";
    tmp(63509) := x"7820";
    tmp(63510) := x"8020";
    tmp(63511) := x"8820";
    tmp(63512) := x"8820";
    tmp(63513) := x"7820";
    tmp(63514) := x"8020";
    tmp(63515) := x"8820";
    tmp(63516) := x"8820";
    tmp(63517) := x"9020";
    tmp(63518) := x"a020";
    tmp(63519) := x"9020";
    tmp(63520) := x"9020";
    tmp(63521) := x"8020";
    tmp(63522) := x"8020";
    tmp(63523) := x"8020";
    tmp(63524) := x"b061";
    tmp(63525) := x"a840";
    tmp(63526) := x"8020";
    tmp(63527) := x"7000";
    tmp(63528) := x"6800";
    tmp(63529) := x"7800";
    tmp(63530) := x"8020";
    tmp(63531) := x"8820";
    tmp(63532) := x"8000";
    tmp(63533) := x"8000";
    tmp(63534) := x"8820";
    tmp(63535) := x"8800";
    tmp(63536) := x"7800";
    tmp(63537) := x"7820";
    tmp(63538) := x"3841";
    tmp(63539) := x"1041";
    tmp(63540) := x"0861";
    tmp(63541) := x"0861";
    tmp(63542) := x"0841";
    tmp(63543) := x"0861";
    tmp(63544) := x"0861";
    tmp(63545) := x"0861";
    tmp(63546) := x"0861";
    tmp(63547) := x"0861";
    tmp(63548) := x"0861";
    tmp(63549) := x"0861";
    tmp(63550) := x"1061";
    tmp(63551) := x"1061";
    tmp(63552) := x"1081";
    tmp(63553) := x"1082";
    tmp(63554) := x"10a2";
    tmp(63555) := x"10a2";
    tmp(63556) := x"18c2";
    tmp(63557) := x"18c3";
    tmp(63558) := x"18e3";
    tmp(63559) := x"20e4";
    tmp(63560) := x"2104";
    tmp(63561) := x"2104";
    tmp(63562) := x"2924";
    tmp(63563) := x"2104";
    tmp(63564) := x"2104";
    tmp(63565) := x"2125";
    tmp(63566) := x"2925";
    tmp(63567) := x"2945";
    tmp(63568) := x"3166";
    tmp(63569) := x"3186";
    tmp(63570) := x"31a7";
    tmp(63571) := x"39c8";
    tmp(63572) := x"39e8";
    tmp(63573) := x"4209";
    tmp(63574) := x"4a2a";
    tmp(63575) := x"4a4a";
    tmp(63576) := x"526b";
    tmp(63577) := x"5a8c";
    tmp(63578) := x"5acd";
    tmp(63579) := x"62cf";
    tmp(63580) := x"6b10";
    tmp(63581) := x"6b50";
    tmp(63582) := x"7391";
    tmp(63583) := x"7bd2";
    tmp(63584) := x"83d3";
    tmp(63585) := x"83f4";
    tmp(63586) := x"8c16";
    tmp(63587) := x"9477";
    tmp(63588) := x"9477";
    tmp(63589) := x"9498";
    tmp(63590) := x"9497";
    tmp(63591) := x"9476";
    tmp(63592) := x"8c55";
    tmp(63593) := x"7c13";
    tmp(63594) := x"7bf2";
    tmp(63595) := x"7bd2";
    tmp(63596) := x"73b1";
    tmp(63597) := x"6b91";
    tmp(63598) := x"6b91";
    tmp(63599) := x"634f";
    tmp(63600) := x"0000";
    tmp(63601) := x"0800";
    tmp(63602) := x"0800";
    tmp(63603) := x"0800";
    tmp(63604) := x"0800";
    tmp(63605) := x"0800";
    tmp(63606) := x"0800";
    tmp(63607) := x"1000";
    tmp(63608) := x"1000";
    tmp(63609) := x"1000";
    tmp(63610) := x"1000";
    tmp(63611) := x"1000";
    tmp(63612) := x"1000";
    tmp(63613) := x"1000";
    tmp(63614) := x"1000";
    tmp(63615) := x"1000";
    tmp(63616) := x"1000";
    tmp(63617) := x"1000";
    tmp(63618) := x"1000";
    tmp(63619) := x"1000";
    tmp(63620) := x"1000";
    tmp(63621) := x"1800";
    tmp(63622) := x"1000";
    tmp(63623) := x"1000";
    tmp(63624) := x"1000";
    tmp(63625) := x"1000";
    tmp(63626) := x"1000";
    tmp(63627) := x"1000";
    tmp(63628) := x"1000";
    tmp(63629) := x"1000";
    tmp(63630) := x"1800";
    tmp(63631) := x"1800";
    tmp(63632) := x"1800";
    tmp(63633) := x"1800";
    tmp(63634) := x"1800";
    tmp(63635) := x"1800";
    tmp(63636) := x"1800";
    tmp(63637) := x"1800";
    tmp(63638) := x"1800";
    tmp(63639) := x"1800";
    tmp(63640) := x"2000";
    tmp(63641) := x"2000";
    tmp(63642) := x"2000";
    tmp(63643) := x"2000";
    tmp(63644) := x"2800";
    tmp(63645) := x"2800";
    tmp(63646) := x"2800";
    tmp(63647) := x"2800";
    tmp(63648) := x"2800";
    tmp(63649) := x"2800";
    tmp(63650) := x"2000";
    tmp(63651) := x"2000";
    tmp(63652) := x"2800";
    tmp(63653) := x"2800";
    tmp(63654) := x"2000";
    tmp(63655) := x"2800";
    tmp(63656) := x"2800";
    tmp(63657) := x"2800";
    tmp(63658) := x"2800";
    tmp(63659) := x"2800";
    tmp(63660) := x"2800";
    tmp(63661) := x"2800";
    tmp(63662) := x"2800";
    tmp(63663) := x"2800";
    tmp(63664) := x"2800";
    tmp(63665) := x"2800";
    tmp(63666) := x"2800";
    tmp(63667) := x"2800";
    tmp(63668) := x"2800";
    tmp(63669) := x"2000";
    tmp(63670) := x"2000";
    tmp(63671) := x"1800";
    tmp(63672) := x"1800";
    tmp(63673) := x"1000";
    tmp(63674) := x"1000";
    tmp(63675) := x"0800";
    tmp(63676) := x"1000";
    tmp(63677) := x"1000";
    tmp(63678) := x"1000";
    tmp(63679) := x"1000";
    tmp(63680) := x"1000";
    tmp(63681) := x"1000";
    tmp(63682) := x"1000";
    tmp(63683) := x"1020";
    tmp(63684) := x"1020";
    tmp(63685) := x"1020";
    tmp(63686) := x"0820";
    tmp(63687) := x"0820";
    tmp(63688) := x"0800";
    tmp(63689) := x"0800";
    tmp(63690) := x"0800";
    tmp(63691) := x"0800";
    tmp(63692) := x"0800";
    tmp(63693) := x"0800";
    tmp(63694) := x"0800";
    tmp(63695) := x"1000";
    tmp(63696) := x"1000";
    tmp(63697) := x"1000";
    tmp(63698) := x"1800";
    tmp(63699) := x"1800";
    tmp(63700) := x"1800";
    tmp(63701) := x"1800";
    tmp(63702) := x"1000";
    tmp(63703) := x"1800";
    tmp(63704) := x"2000";
    tmp(63705) := x"2000";
    tmp(63706) := x"1800";
    tmp(63707) := x"1000";
    tmp(63708) := x"0800";
    tmp(63709) := x"0800";
    tmp(63710) := x"1800";
    tmp(63711) := x"2000";
    tmp(63712) := x"2800";
    tmp(63713) := x"2800";
    tmp(63714) := x"2000";
    tmp(63715) := x"2800";
    tmp(63716) := x"3000";
    tmp(63717) := x"3000";
    tmp(63718) := x"3000";
    tmp(63719) := x"4000";
    tmp(63720) := x"4000";
    tmp(63721) := x"4000";
    tmp(63722) := x"5000";
    tmp(63723) := x"5800";
    tmp(63724) := x"6000";
    tmp(63725) := x"6000";
    tmp(63726) := x"5800";
    tmp(63727) := x"5000";
    tmp(63728) := x"6000";
    tmp(63729) := x"5800";
    tmp(63730) := x"5800";
    tmp(63731) := x"6000";
    tmp(63732) := x"5800";
    tmp(63733) := x"5800";
    tmp(63734) := x"6000";
    tmp(63735) := x"6000";
    tmp(63736) := x"6000";
    tmp(63737) := x"7000";
    tmp(63738) := x"7000";
    tmp(63739) := x"7000";
    tmp(63740) := x"6800";
    tmp(63741) := x"5800";
    tmp(63742) := x"6000";
    tmp(63743) := x"6820";
    tmp(63744) := x"6000";
    tmp(63745) := x"6800";
    tmp(63746) := x"6000";
    tmp(63747) := x"7020";
    tmp(63748) := x"8820";
    tmp(63749) := x"7820";
    tmp(63750) := x"7820";
    tmp(63751) := x"7820";
    tmp(63752) := x"7820";
    tmp(63753) := x"7020";
    tmp(63754) := x"7820";
    tmp(63755) := x"9020";
    tmp(63756) := x"8820";
    tmp(63757) := x"9020";
    tmp(63758) := x"a020";
    tmp(63759) := x"a040";
    tmp(63760) := x"a040";
    tmp(63761) := x"8820";
    tmp(63762) := x"7800";
    tmp(63763) := x"7020";
    tmp(63764) := x"9020";
    tmp(63765) := x"8820";
    tmp(63766) := x"8820";
    tmp(63767) := x"6800";
    tmp(63768) := x"7000";
    tmp(63769) := x"7800";
    tmp(63770) := x"7000";
    tmp(63771) := x"7800";
    tmp(63772) := x"8020";
    tmp(63773) := x"8020";
    tmp(63774) := x"8820";
    tmp(63775) := x"8020";
    tmp(63776) := x"7820";
    tmp(63777) := x"5040";
    tmp(63778) := x"1841";
    tmp(63779) := x"1041";
    tmp(63780) := x"0861";
    tmp(63781) := x"0841";
    tmp(63782) := x"0841";
    tmp(63783) := x"0861";
    tmp(63784) := x"0861";
    tmp(63785) := x"0861";
    tmp(63786) := x"0861";
    tmp(63787) := x"0861";
    tmp(63788) := x"1061";
    tmp(63789) := x"1081";
    tmp(63790) := x"1081";
    tmp(63791) := x"1082";
    tmp(63792) := x"10a2";
    tmp(63793) := x"10a2";
    tmp(63794) := x"18a2";
    tmp(63795) := x"18c3";
    tmp(63796) := x"18e3";
    tmp(63797) := x"20e4";
    tmp(63798) := x"2104";
    tmp(63799) := x"2925";
    tmp(63800) := x"2925";
    tmp(63801) := x"2945";
    tmp(63802) := x"2945";
    tmp(63803) := x"2945";
    tmp(63804) := x"2945";
    tmp(63805) := x"2945";
    tmp(63806) := x"2966";
    tmp(63807) := x"3166";
    tmp(63808) := x"39a7";
    tmp(63809) := x"39a7";
    tmp(63810) := x"39e8";
    tmp(63811) := x"4209";
    tmp(63812) := x"4a2a";
    tmp(63813) := x"524b";
    tmp(63814) := x"524b";
    tmp(63815) := x"528c";
    tmp(63816) := x"5acd";
    tmp(63817) := x"62ee";
    tmp(63818) := x"6aef";
    tmp(63819) := x"7350";
    tmp(63820) := x"7b72";
    tmp(63821) := x"7b92";
    tmp(63822) := x"83d3";
    tmp(63823) := x"8c15";
    tmp(63824) := x"9456";
    tmp(63825) := x"9477";
    tmp(63826) := x"9497";
    tmp(63827) := x"9cd8";
    tmp(63828) := x"9cd8";
    tmp(63829) := x"a53a";
    tmp(63830) := x"9cf9";
    tmp(63831) := x"9cd8";
    tmp(63832) := x"9497";
    tmp(63833) := x"8c75";
    tmp(63834) := x"8c54";
    tmp(63835) := x"8c33";
    tmp(63836) := x"7bb2";
    tmp(63837) := x"73d2";
    tmp(63838) := x"6b91";
    tmp(63839) := x"6b6f";
    tmp(63840) := x"0000";
    tmp(63841) := x"0800";
    tmp(63842) := x"0800";
    tmp(63843) := x"0800";
    tmp(63844) := x"0800";
    tmp(63845) := x"0800";
    tmp(63846) := x"1000";
    tmp(63847) := x"1000";
    tmp(63848) := x"1000";
    tmp(63849) := x"1000";
    tmp(63850) := x"1000";
    tmp(63851) := x"1000";
    tmp(63852) := x"1000";
    tmp(63853) := x"1000";
    tmp(63854) := x"1000";
    tmp(63855) := x"1000";
    tmp(63856) := x"1000";
    tmp(63857) := x"1000";
    tmp(63858) := x"1000";
    tmp(63859) := x"1000";
    tmp(63860) := x"1000";
    tmp(63861) := x"1800";
    tmp(63862) := x"1800";
    tmp(63863) := x"1800";
    tmp(63864) := x"1000";
    tmp(63865) := x"1000";
    tmp(63866) := x"1000";
    tmp(63867) := x"1000";
    tmp(63868) := x"1000";
    tmp(63869) := x"1000";
    tmp(63870) := x"1800";
    tmp(63871) := x"1800";
    tmp(63872) := x"1800";
    tmp(63873) := x"1800";
    tmp(63874) := x"1800";
    tmp(63875) := x"1800";
    tmp(63876) := x"1000";
    tmp(63877) := x"1800";
    tmp(63878) := x"1800";
    tmp(63879) := x"1800";
    tmp(63880) := x"1800";
    tmp(63881) := x"1800";
    tmp(63882) := x"2000";
    tmp(63883) := x"2000";
    tmp(63884) := x"2000";
    tmp(63885) := x"2000";
    tmp(63886) := x"2800";
    tmp(63887) := x"2800";
    tmp(63888) := x"2800";
    tmp(63889) := x"2800";
    tmp(63890) := x"2800";
    tmp(63891) := x"2000";
    tmp(63892) := x"2000";
    tmp(63893) := x"2000";
    tmp(63894) := x"2000";
    tmp(63895) := x"2000";
    tmp(63896) := x"2000";
    tmp(63897) := x"2800";
    tmp(63898) := x"2800";
    tmp(63899) := x"2800";
    tmp(63900) := x"2000";
    tmp(63901) := x"2000";
    tmp(63902) := x"2800";
    tmp(63903) := x"2000";
    tmp(63904) := x"2800";
    tmp(63905) := x"2800";
    tmp(63906) := x"2800";
    tmp(63907) := x"2800";
    tmp(63908) := x"2800";
    tmp(63909) := x"2800";
    tmp(63910) := x"2000";
    tmp(63911) := x"1800";
    tmp(63912) := x"1000";
    tmp(63913) := x"1000";
    tmp(63914) := x"1000";
    tmp(63915) := x"1800";
    tmp(63916) := x"1000";
    tmp(63917) := x"1000";
    tmp(63918) := x"1000";
    tmp(63919) := x"1000";
    tmp(63920) := x"1000";
    tmp(63921) := x"1000";
    tmp(63922) := x"1000";
    tmp(63923) := x"1000";
    tmp(63924) := x"1020";
    tmp(63925) := x"0820";
    tmp(63926) := x"0820";
    tmp(63927) := x"0820";
    tmp(63928) := x"0800";
    tmp(63929) := x"0800";
    tmp(63930) := x"0800";
    tmp(63931) := x"0800";
    tmp(63932) := x"0800";
    tmp(63933) := x"0800";
    tmp(63934) := x"1000";
    tmp(63935) := x"1000";
    tmp(63936) := x"1800";
    tmp(63937) := x"1800";
    tmp(63938) := x"1800";
    tmp(63939) := x"1800";
    tmp(63940) := x"1800";
    tmp(63941) := x"1800";
    tmp(63942) := x"1800";
    tmp(63943) := x"1800";
    tmp(63944) := x"1800";
    tmp(63945) := x"1800";
    tmp(63946) := x"1000";
    tmp(63947) := x"0800";
    tmp(63948) := x"0800";
    tmp(63949) := x"1000";
    tmp(63950) := x"1800";
    tmp(63951) := x"2000";
    tmp(63952) := x"2000";
    tmp(63953) := x"2000";
    tmp(63954) := x"2000";
    tmp(63955) := x"2800";
    tmp(63956) := x"2800";
    tmp(63957) := x"3000";
    tmp(63958) := x"3000";
    tmp(63959) := x"3800";
    tmp(63960) := x"4000";
    tmp(63961) := x"4000";
    tmp(63962) := x"4800";
    tmp(63963) := x"5800";
    tmp(63964) := x"5800";
    tmp(63965) := x"5800";
    tmp(63966) := x"5000";
    tmp(63967) := x"5800";
    tmp(63968) := x"6000";
    tmp(63969) := x"5800";
    tmp(63970) := x"5000";
    tmp(63971) := x"5800";
    tmp(63972) := x"5000";
    tmp(63973) := x"5800";
    tmp(63974) := x"5800";
    tmp(63975) := x"6000";
    tmp(63976) := x"6000";
    tmp(63977) := x"7800";
    tmp(63978) := x"6800";
    tmp(63979) := x"7000";
    tmp(63980) := x"6000";
    tmp(63981) := x"5800";
    tmp(63982) := x"6000";
    tmp(63983) := x"6820";
    tmp(63984) := x"6800";
    tmp(63985) := x"7000";
    tmp(63986) := x"6800";
    tmp(63987) := x"8020";
    tmp(63988) := x"8820";
    tmp(63989) := x"8020";
    tmp(63990) := x"7000";
    tmp(63991) := x"7020";
    tmp(63992) := x"7820";
    tmp(63993) := x"6800";
    tmp(63994) := x"8820";
    tmp(63995) := x"8820";
    tmp(63996) := x"8820";
    tmp(63997) := x"9020";
    tmp(63998) := x"a840";
    tmp(63999) := x"b861";
    tmp(64000) := x"b061";
    tmp(64001) := x"8820";
    tmp(64002) := x"7820";
    tmp(64003) := x"7820";
    tmp(64004) := x"9020";
    tmp(64005) := x"9820";
    tmp(64006) := x"8020";
    tmp(64007) := x"7820";
    tmp(64008) := x"7000";
    tmp(64009) := x"7800";
    tmp(64010) := x"6800";
    tmp(64011) := x"7800";
    tmp(64012) := x"8820";
    tmp(64013) := x"8820";
    tmp(64014) := x"9820";
    tmp(64015) := x"7020";
    tmp(64016) := x"3840";
    tmp(64017) := x"2041";
    tmp(64018) := x"1041";
    tmp(64019) := x"0841";
    tmp(64020) := x"0841";
    tmp(64021) := x"0841";
    tmp(64022) := x"0841";
    tmp(64023) := x"0861";
    tmp(64024) := x"1061";
    tmp(64025) := x"1061";
    tmp(64026) := x"1061";
    tmp(64027) := x"1081";
    tmp(64028) := x"1082";
    tmp(64029) := x"1082";
    tmp(64030) := x"10a2";
    tmp(64031) := x"10a2";
    tmp(64032) := x"18c2";
    tmp(64033) := x"18c3";
    tmp(64034) := x"18e3";
    tmp(64035) := x"2104";
    tmp(64036) := x"2104";
    tmp(64037) := x"2925";
    tmp(64038) := x"2945";
    tmp(64039) := x"2946";
    tmp(64040) := x"3166";
    tmp(64041) := x"3166";
    tmp(64042) := x"3166";
    tmp(64043) := x"3166";
    tmp(64044) := x"3166";
    tmp(64045) := x"3187";
    tmp(64046) := x"3187";
    tmp(64047) := x"39a7";
    tmp(64048) := x"39c8";
    tmp(64049) := x"4209";
    tmp(64050) := x"4a4a";
    tmp(64051) := x"4a4b";
    tmp(64052) := x"524b";
    tmp(64053) := x"526c";
    tmp(64054) := x"5a8d";
    tmp(64055) := x"62ce";
    tmp(64056) := x"6b2f";
    tmp(64057) := x"7351";
    tmp(64058) := x"7b92";
    tmp(64059) := x"83b3";
    tmp(64060) := x"83b4";
    tmp(64061) := x"8c16";
    tmp(64062) := x"9456";
    tmp(64063) := x"9477";
    tmp(64064) := x"9c98";
    tmp(64065) := x"a4d9";
    tmp(64066) := x"ad3b";
    tmp(64067) := x"b57c";
    tmp(64068) := x"a53b";
    tmp(64069) := x"b59d";
    tmp(64070) := x"a55b";
    tmp(64071) := x"a53a";
    tmp(64072) := x"94f8";
    tmp(64073) := x"94b7";
    tmp(64074) := x"9496";
    tmp(64075) := x"8c54";
    tmp(64076) := x"8413";
    tmp(64077) := x"73b1";
    tmp(64078) := x"6b91";
    tmp(64079) := x"6bb1";
    tmp(64080) := x"0000";
    tmp(64081) := x"0800";
    tmp(64082) := x"0800";
    tmp(64083) := x"0800";
    tmp(64084) := x"0800";
    tmp(64085) := x"1000";
    tmp(64086) := x"1000";
    tmp(64087) := x"0800";
    tmp(64088) := x"1000";
    tmp(64089) := x"1000";
    tmp(64090) := x"1000";
    tmp(64091) := x"1000";
    tmp(64092) := x"1000";
    tmp(64093) := x"1000";
    tmp(64094) := x"1000";
    tmp(64095) := x"1000";
    tmp(64096) := x"1000";
    tmp(64097) := x"1000";
    tmp(64098) := x"1000";
    tmp(64099) := x"1000";
    tmp(64100) := x"1000";
    tmp(64101) := x"1800";
    tmp(64102) := x"1800";
    tmp(64103) := x"1800";
    tmp(64104) := x"1800";
    tmp(64105) := x"1000";
    tmp(64106) := x"1000";
    tmp(64107) := x"1000";
    tmp(64108) := x"1000";
    tmp(64109) := x"1000";
    tmp(64110) := x"1000";
    tmp(64111) := x"1800";
    tmp(64112) := x"1800";
    tmp(64113) := x"1800";
    tmp(64114) := x"1800";
    tmp(64115) := x"1800";
    tmp(64116) := x"1800";
    tmp(64117) := x"1800";
    tmp(64118) := x"1800";
    tmp(64119) := x"1800";
    tmp(64120) := x"1800";
    tmp(64121) := x"2000";
    tmp(64122) := x"2000";
    tmp(64123) := x"2000";
    tmp(64124) := x"2000";
    tmp(64125) := x"2000";
    tmp(64126) := x"2000";
    tmp(64127) := x"2000";
    tmp(64128) := x"2000";
    tmp(64129) := x"2000";
    tmp(64130) := x"2000";
    tmp(64131) := x"2000";
    tmp(64132) := x"2000";
    tmp(64133) := x"2000";
    tmp(64134) := x"2000";
    tmp(64135) := x"2000";
    tmp(64136) := x"2000";
    tmp(64137) := x"2000";
    tmp(64138) := x"2000";
    tmp(64139) := x"2000";
    tmp(64140) := x"2000";
    tmp(64141) := x"2000";
    tmp(64142) := x"2000";
    tmp(64143) := x"2000";
    tmp(64144) := x"2000";
    tmp(64145) := x"2000";
    tmp(64146) := x"2000";
    tmp(64147) := x"2000";
    tmp(64148) := x"2000";
    tmp(64149) := x"2000";
    tmp(64150) := x"2000";
    tmp(64151) := x"1800";
    tmp(64152) := x"1000";
    tmp(64153) := x"1000";
    tmp(64154) := x"1800";
    tmp(64155) := x"1800";
    tmp(64156) := x"1000";
    tmp(64157) := x"1000";
    tmp(64158) := x"1000";
    tmp(64159) := x"1000";
    tmp(64160) := x"1000";
    tmp(64161) := x"1000";
    tmp(64162) := x"1000";
    tmp(64163) := x"1020";
    tmp(64164) := x"0820";
    tmp(64165) := x"0820";
    tmp(64166) := x"0800";
    tmp(64167) := x"0820";
    tmp(64168) := x"0800";
    tmp(64169) := x"0800";
    tmp(64170) := x"0800";
    tmp(64171) := x"0800";
    tmp(64172) := x"0800";
    tmp(64173) := x"1000";
    tmp(64174) := x"1000";
    tmp(64175) := x"1000";
    tmp(64176) := x"1800";
    tmp(64177) := x"1800";
    tmp(64178) := x"2000";
    tmp(64179) := x"2000";
    tmp(64180) := x"1800";
    tmp(64181) := x"1800";
    tmp(64182) := x"1800";
    tmp(64183) := x"1800";
    tmp(64184) := x"1800";
    tmp(64185) := x"1000";
    tmp(64186) := x"0800";
    tmp(64187) := x"0800";
    tmp(64188) := x"0800";
    tmp(64189) := x"1000";
    tmp(64190) := x"1800";
    tmp(64191) := x"2000";
    tmp(64192) := x"2000";
    tmp(64193) := x"2800";
    tmp(64194) := x"2800";
    tmp(64195) := x"2800";
    tmp(64196) := x"3000";
    tmp(64197) := x"3000";
    tmp(64198) := x"3000";
    tmp(64199) := x"3800";
    tmp(64200) := x"4000";
    tmp(64201) := x"3800";
    tmp(64202) := x"4800";
    tmp(64203) := x"5800";
    tmp(64204) := x"6000";
    tmp(64205) := x"5800";
    tmp(64206) := x"5000";
    tmp(64207) := x"5800";
    tmp(64208) := x"5800";
    tmp(64209) := x"5800";
    tmp(64210) := x"5800";
    tmp(64211) := x"5000";
    tmp(64212) := x"5800";
    tmp(64213) := x"5800";
    tmp(64214) := x"6000";
    tmp(64215) := x"6000";
    tmp(64216) := x"6800";
    tmp(64217) := x"6800";
    tmp(64218) := x"7000";
    tmp(64219) := x"7000";
    tmp(64220) := x"6000";
    tmp(64221) := x"5800";
    tmp(64222) := x"6800";
    tmp(64223) := x"7020";
    tmp(64224) := x"7020";
    tmp(64225) := x"7020";
    tmp(64226) := x"7020";
    tmp(64227) := x"8020";
    tmp(64228) := x"7820";
    tmp(64229) := x"7020";
    tmp(64230) := x"5800";
    tmp(64231) := x"8020";
    tmp(64232) := x"6800";
    tmp(64233) := x"7820";
    tmp(64234) := x"8820";
    tmp(64235) := x"8820";
    tmp(64236) := x"9020";
    tmp(64237) := x"a020";
    tmp(64238) := x"a840";
    tmp(64239) := x"b040";
    tmp(64240) := x"b041";
    tmp(64241) := x"8020";
    tmp(64242) := x"8020";
    tmp(64243) := x"8020";
    tmp(64244) := x"7800";
    tmp(64245) := x"8800";
    tmp(64246) := x"8020";
    tmp(64247) := x"8820";
    tmp(64248) := x"7800";
    tmp(64249) := x"7000";
    tmp(64250) := x"6000";
    tmp(64251) := x"7800";
    tmp(64252) := x"8820";
    tmp(64253) := x"8820";
    tmp(64254) := x"9020";
    tmp(64255) := x"3840";
    tmp(64256) := x"1040";
    tmp(64257) := x"1041";
    tmp(64258) := x"0841";
    tmp(64259) := x"0841";
    tmp(64260) := x"0861";
    tmp(64261) := x"0861";
    tmp(64262) := x"1061";
    tmp(64263) := x"1061";
    tmp(64264) := x"1061";
    tmp(64265) := x"1082";
    tmp(64266) := x"1082";
    tmp(64267) := x"1082";
    tmp(64268) := x"10a2";
    tmp(64269) := x"18a2";
    tmp(64270) := x"18a2";
    tmp(64271) := x"18c3";
    tmp(64272) := x"18c3";
    tmp(64273) := x"2104";
    tmp(64274) := x"2104";
    tmp(64275) := x"2925";
    tmp(64276) := x"2945";
    tmp(64277) := x"2966";
    tmp(64278) := x"3166";
    tmp(64279) := x"3187";
    tmp(64280) := x"3187";
    tmp(64281) := x"31a7";
    tmp(64282) := x"31a7";
    tmp(64283) := x"39a7";
    tmp(64284) := x"39a7";
    tmp(64285) := x"39a8";
    tmp(64286) := x"39c8";
    tmp(64287) := x"41e9";
    tmp(64288) := x"4a2a";
    tmp(64289) := x"4a2a";
    tmp(64290) := x"526b";
    tmp(64291) := x"526c";
    tmp(64292) := x"5aad";
    tmp(64293) := x"62cd";
    tmp(64294) := x"6aef";
    tmp(64295) := x"7331";
    tmp(64296) := x"7b72";
    tmp(64297) := x"83d3";
    tmp(64298) := x"8bf5";
    tmp(64299) := x"8bf5";
    tmp(64300) := x"9457";
    tmp(64301) := x"9c98";
    tmp(64302) := x"a4f9";
    tmp(64303) := x"a4fa";
    tmp(64304) := x"ad3d";
    tmp(64305) := x"b55d";
    tmp(64306) := x"bdde";
    tmp(64307) := x"bdbd";
    tmp(64308) := x"bdde";
    tmp(64309) := x"b5bd";
    tmp(64310) := x"bddd";
    tmp(64311) := x"ad7b";
    tmp(64312) := x"9d19";
    tmp(64313) := x"9cd7";
    tmp(64314) := x"9496";
    tmp(64315) := x"8c54";
    tmp(64316) := x"7bf3";
    tmp(64317) := x"73d2";
    tmp(64318) := x"73d2";
    tmp(64319) := x"7392";
    tmp(64320) := x"0000";
    tmp(64321) := x"0800";
    tmp(64322) := x"0800";
    tmp(64323) := x"0800";
    tmp(64324) := x"0800";
    tmp(64325) := x"0800";
    tmp(64326) := x"0800";
    tmp(64327) := x"0800";
    tmp(64328) := x"1000";
    tmp(64329) := x"1000";
    tmp(64330) := x"1000";
    tmp(64331) := x"1000";
    tmp(64332) := x"1000";
    tmp(64333) := x"1000";
    tmp(64334) := x"1000";
    tmp(64335) := x"1000";
    tmp(64336) := x"1000";
    tmp(64337) := x"1000";
    tmp(64338) := x"1000";
    tmp(64339) := x"1000";
    tmp(64340) := x"1800";
    tmp(64341) := x"1800";
    tmp(64342) := x"1800";
    tmp(64343) := x"1800";
    tmp(64344) := x"2000";
    tmp(64345) := x"1800";
    tmp(64346) := x"1000";
    tmp(64347) := x"1000";
    tmp(64348) := x"1000";
    tmp(64349) := x"1000";
    tmp(64350) := x"1800";
    tmp(64351) := x"1800";
    tmp(64352) := x"1800";
    tmp(64353) := x"1800";
    tmp(64354) := x"1800";
    tmp(64355) := x"1800";
    tmp(64356) := x"1800";
    tmp(64357) := x"1800";
    tmp(64358) := x"1800";
    tmp(64359) := x"1800";
    tmp(64360) := x"1800";
    tmp(64361) := x"1800";
    tmp(64362) := x"1800";
    tmp(64363) := x"1800";
    tmp(64364) := x"2000";
    tmp(64365) := x"2000";
    tmp(64366) := x"2000";
    tmp(64367) := x"2000";
    tmp(64368) := x"2000";
    tmp(64369) := x"2000";
    tmp(64370) := x"2000";
    tmp(64371) := x"2000";
    tmp(64372) := x"2000";
    tmp(64373) := x"2000";
    tmp(64374) := x"2000";
    tmp(64375) := x"1800";
    tmp(64376) := x"1800";
    tmp(64377) := x"1800";
    tmp(64378) := x"1800";
    tmp(64379) := x"1800";
    tmp(64380) := x"2000";
    tmp(64381) := x"2000";
    tmp(64382) := x"2000";
    tmp(64383) := x"2000";
    tmp(64384) := x"2000";
    tmp(64385) := x"2000";
    tmp(64386) := x"2000";
    tmp(64387) := x"2000";
    tmp(64388) := x"2000";
    tmp(64389) := x"2000";
    tmp(64390) := x"1800";
    tmp(64391) := x"1800";
    tmp(64392) := x"1800";
    tmp(64393) := x"1800";
    tmp(64394) := x"1800";
    tmp(64395) := x"1800";
    tmp(64396) := x"1000";
    tmp(64397) := x"1000";
    tmp(64398) := x"1000";
    tmp(64399) := x"1000";
    tmp(64400) := x"1000";
    tmp(64401) := x"1000";
    tmp(64402) := x"0800";
    tmp(64403) := x"0800";
    tmp(64404) := x"0820";
    tmp(64405) := x"0800";
    tmp(64406) := x"0800";
    tmp(64407) := x"0800";
    tmp(64408) := x"0800";
    tmp(64409) := x"0800";
    tmp(64410) := x"0800";
    tmp(64411) := x"0800";
    tmp(64412) := x"1000";
    tmp(64413) := x"1000";
    tmp(64414) := x"1000";
    tmp(64415) := x"1000";
    tmp(64416) := x"1000";
    tmp(64417) := x"1000";
    tmp(64418) := x"1800";
    tmp(64419) := x"1800";
    tmp(64420) := x"1800";
    tmp(64421) := x"1800";
    tmp(64422) := x"1000";
    tmp(64423) := x"1000";
    tmp(64424) := x"0800";
    tmp(64425) := x"0800";
    tmp(64426) := x"0800";
    tmp(64427) := x"0800";
    tmp(64428) := x"0800";
    tmp(64429) := x"0800";
    tmp(64430) := x"1000";
    tmp(64431) := x"2000";
    tmp(64432) := x"2800";
    tmp(64433) := x"2800";
    tmp(64434) := x"2000";
    tmp(64435) := x"2000";
    tmp(64436) := x"3000";
    tmp(64437) := x"3800";
    tmp(64438) := x"3800";
    tmp(64439) := x"4000";
    tmp(64440) := x"3800";
    tmp(64441) := x"3800";
    tmp(64442) := x"4800";
    tmp(64443) := x"5800";
    tmp(64444) := x"5800";
    tmp(64445) := x"5000";
    tmp(64446) := x"5000";
    tmp(64447) := x"5800";
    tmp(64448) := x"5800";
    tmp(64449) := x"5000";
    tmp(64450) := x"5000";
    tmp(64451) := x"5800";
    tmp(64452) := x"5800";
    tmp(64453) := x"5800";
    tmp(64454) := x"5800";
    tmp(64455) := x"5800";
    tmp(64456) := x"6800";
    tmp(64457) := x"6000";
    tmp(64458) := x"7000";
    tmp(64459) := x"6800";
    tmp(64460) := x"5800";
    tmp(64461) := x"5800";
    tmp(64462) := x"6800";
    tmp(64463) := x"7020";
    tmp(64464) := x"7820";
    tmp(64465) := x"7820";
    tmp(64466) := x"7820";
    tmp(64467) := x"7020";
    tmp(64468) := x"6820";
    tmp(64469) := x"7020";
    tmp(64470) := x"5000";
    tmp(64471) := x"6000";
    tmp(64472) := x"7020";
    tmp(64473) := x"8020";
    tmp(64474) := x"8020";
    tmp(64475) := x"9020";
    tmp(64476) := x"a020";
    tmp(64477) := x"a820";
    tmp(64478) := x"b040";
    tmp(64479) := x"9840";
    tmp(64480) := x"a861";
    tmp(64481) := x"7820";
    tmp(64482) := x"8820";
    tmp(64483) := x"7000";
    tmp(64484) := x"7000";
    tmp(64485) := x"7000";
    tmp(64486) := x"8020";
    tmp(64487) := x"8820";
    tmp(64488) := x"8020";
    tmp(64489) := x"7000";
    tmp(64490) := x"7000";
    tmp(64491) := x"7820";
    tmp(64492) := x"8020";
    tmp(64493) := x"7820";
    tmp(64494) := x"5040";
    tmp(64495) := x"1840";
    tmp(64496) := x"0840";
    tmp(64497) := x"0841";
    tmp(64498) := x"0841";
    tmp(64499) := x"0841";
    tmp(64500) := x"0861";
    tmp(64501) := x"1061";
    tmp(64502) := x"1061";
    tmp(64503) := x"1081";
    tmp(64504) := x"1082";
    tmp(64505) := x"10a2";
    tmp(64506) := x"10a2";
    tmp(64507) := x"18a2";
    tmp(64508) := x"18a2";
    tmp(64509) := x"18c3";
    tmp(64510) := x"18e3";
    tmp(64511) := x"20e3";
    tmp(64512) := x"2104";
    tmp(64513) := x"2124";
    tmp(64514) := x"2925";
    tmp(64515) := x"2946";
    tmp(64516) := x"3166";
    tmp(64517) := x"3187";
    tmp(64518) := x"39a7";
    tmp(64519) := x"39a7";
    tmp(64520) := x"39a8";
    tmp(64521) := x"39c8";
    tmp(64522) := x"39c8";
    tmp(64523) := x"39c8";
    tmp(64524) := x"39c9";
    tmp(64525) := x"41e9";
    tmp(64526) := x"4a09";
    tmp(64527) := x"4a2a";
    tmp(64528) := x"526b";
    tmp(64529) := x"5a8c";
    tmp(64530) := x"5aad";
    tmp(64531) := x"62ce";
    tmp(64532) := x"6b0f";
    tmp(64533) := x"7350";
    tmp(64534) := x"7b91";
    tmp(64535) := x"83b3";
    tmp(64536) := x"8bf4";
    tmp(64537) := x"8c15";
    tmp(64538) := x"9457";
    tmp(64539) := x"9c78";
    tmp(64540) := x"acfb";
    tmp(64541) := x"b55d";
    tmp(64542) := x"b57d";
    tmp(64543) := x"bd7d";
    tmp(64544) := x"bdbd";
    tmp(64545) := x"c5ff";
    tmp(64546) := x"c5ff";
    tmp(64547) := x"c61f";
    tmp(64548) := x"c5ff";
    tmp(64549) := x"bdff";
    tmp(64550) := x"b5be";
    tmp(64551) := x"b59d";
    tmp(64552) := x"ad5b";
    tmp(64553) := x"9cd7";
    tmp(64554) := x"9476";
    tmp(64555) := x"8c55";
    tmp(64556) := x"7c13";
    tmp(64557) := x"7bf3";
    tmp(64558) := x"73d2";
    tmp(64559) := x"6bb1";
    tmp(64560) := x"0000";
    tmp(64561) := x"0800";
    tmp(64562) := x"0800";
    tmp(64563) := x"0800";
    tmp(64564) := x"0800";
    tmp(64565) := x"0800";
    tmp(64566) := x"0800";
    tmp(64567) := x"1000";
    tmp(64568) := x"1000";
    tmp(64569) := x"1000";
    tmp(64570) := x"1000";
    tmp(64571) := x"1000";
    tmp(64572) := x"1000";
    tmp(64573) := x"1000";
    tmp(64574) := x"1000";
    tmp(64575) := x"1000";
    tmp(64576) := x"1000";
    tmp(64577) := x"1000";
    tmp(64578) := x"1000";
    tmp(64579) := x"1800";
    tmp(64580) := x"1800";
    tmp(64581) := x"1800";
    tmp(64582) := x"1800";
    tmp(64583) := x"1800";
    tmp(64584) := x"1800";
    tmp(64585) := x"1800";
    tmp(64586) := x"1800";
    tmp(64587) := x"1800";
    tmp(64588) := x"1000";
    tmp(64589) := x"1000";
    tmp(64590) := x"1800";
    tmp(64591) := x"1800";
    tmp(64592) := x"1800";
    tmp(64593) := x"1800";
    tmp(64594) := x"1800";
    tmp(64595) := x"1800";
    tmp(64596) := x"1800";
    tmp(64597) := x"1800";
    tmp(64598) := x"1800";
    tmp(64599) := x"1800";
    tmp(64600) := x"1800";
    tmp(64601) := x"1800";
    tmp(64602) := x"1800";
    tmp(64603) := x"1800";
    tmp(64604) := x"1800";
    tmp(64605) := x"2000";
    tmp(64606) := x"2000";
    tmp(64607) := x"2000";
    tmp(64608) := x"2000";
    tmp(64609) := x"2000";
    tmp(64610) := x"2000";
    tmp(64611) := x"2000";
    tmp(64612) := x"2000";
    tmp(64613) := x"2000";
    tmp(64614) := x"2000";
    tmp(64615) := x"1800";
    tmp(64616) := x"1800";
    tmp(64617) := x"1800";
    tmp(64618) := x"1800";
    tmp(64619) := x"1800";
    tmp(64620) := x"1800";
    tmp(64621) := x"1800";
    tmp(64622) := x"2000";
    tmp(64623) := x"2000";
    tmp(64624) := x"1800";
    tmp(64625) := x"1800";
    tmp(64626) := x"2000";
    tmp(64627) := x"1800";
    tmp(64628) := x"1800";
    tmp(64629) := x"1800";
    tmp(64630) := x"1800";
    tmp(64631) := x"1800";
    tmp(64632) := x"1800";
    tmp(64633) := x"1800";
    tmp(64634) := x"1000";
    tmp(64635) := x"1000";
    tmp(64636) := x"0800";
    tmp(64637) := x"0800";
    tmp(64638) := x"0800";
    tmp(64639) := x"0800";
    tmp(64640) := x"0800";
    tmp(64641) := x"0800";
    tmp(64642) := x"0820";
    tmp(64643) := x"0820";
    tmp(64644) := x"0820";
    tmp(64645) := x"0800";
    tmp(64646) := x"0800";
    tmp(64647) := x"0800";
    tmp(64648) := x"0800";
    tmp(64649) := x"0800";
    tmp(64650) := x"0800";
    tmp(64651) := x"0800";
    tmp(64652) := x"1000";
    tmp(64653) := x"1000";
    tmp(64654) := x"1000";
    tmp(64655) := x"1000";
    tmp(64656) := x"1000";
    tmp(64657) := x"1000";
    tmp(64658) := x"1000";
    tmp(64659) := x"1000";
    tmp(64660) := x"1000";
    tmp(64661) := x"1000";
    tmp(64662) := x"1000";
    tmp(64663) := x"1000";
    tmp(64664) := x"1000";
    tmp(64665) := x"1000";
    tmp(64666) := x"1000";
    tmp(64667) := x"0800";
    tmp(64668) := x"0800";
    tmp(64669) := x"0800";
    tmp(64670) := x"1000";
    tmp(64671) := x"1800";
    tmp(64672) := x"1800";
    tmp(64673) := x"2000";
    tmp(64674) := x"2800";
    tmp(64675) := x"3000";
    tmp(64676) := x"3800";
    tmp(64677) := x"3800";
    tmp(64678) := x"3800";
    tmp(64679) := x"3800";
    tmp(64680) := x"3800";
    tmp(64681) := x"4000";
    tmp(64682) := x"4800";
    tmp(64683) := x"5800";
    tmp(64684) := x"5000";
    tmp(64685) := x"5000";
    tmp(64686) := x"5000";
    tmp(64687) := x"5000";
    tmp(64688) := x"5000";
    tmp(64689) := x"5000";
    tmp(64690) := x"5800";
    tmp(64691) := x"5800";
    tmp(64692) := x"5800";
    tmp(64693) := x"5800";
    tmp(64694) := x"5800";
    tmp(64695) := x"6000";
    tmp(64696) := x"6000";
    tmp(64697) := x"6800";
    tmp(64698) := x"7800";
    tmp(64699) := x"6000";
    tmp(64700) := x"5800";
    tmp(64701) := x"6000";
    tmp(64702) := x"6800";
    tmp(64703) := x"6800";
    tmp(64704) := x"7820";
    tmp(64705) := x"7820";
    tmp(64706) := x"7020";
    tmp(64707) := x"6800";
    tmp(64708) := x"5800";
    tmp(64709) := x"6000";
    tmp(64710) := x"5000";
    tmp(64711) := x"5800";
    tmp(64712) := x"7020";
    tmp(64713) := x"8020";
    tmp(64714) := x"8820";
    tmp(64715) := x"a020";
    tmp(64716) := x"b020";
    tmp(64717) := x"c840";
    tmp(64718) := x"b841";
    tmp(64719) := x"8020";
    tmp(64720) := x"7820";
    tmp(64721) := x"8840";
    tmp(64722) := x"7820";
    tmp(64723) := x"6800";
    tmp(64724) := x"6000";
    tmp(64725) := x"6800";
    tmp(64726) := x"9020";
    tmp(64727) := x"9020";
    tmp(64728) := x"8820";
    tmp(64729) := x"7820";
    tmp(64730) := x"8020";
    tmp(64731) := x"8020";
    tmp(64732) := x"8820";
    tmp(64733) := x"5820";
    tmp(64734) := x"1840";
    tmp(64735) := x"0840";
    tmp(64736) := x"0840";
    tmp(64737) := x"0840";
    tmp(64738) := x"0841";
    tmp(64739) := x"0841";
    tmp(64740) := x"0861";
    tmp(64741) := x"1061";
    tmp(64742) := x"1081";
    tmp(64743) := x"1082";
    tmp(64744) := x"10a2";
    tmp(64745) := x"10a2";
    tmp(64746) := x"18c3";
    tmp(64747) := x"18c3";
    tmp(64748) := x"18c3";
    tmp(64749) := x"20e3";
    tmp(64750) := x"20e4";
    tmp(64751) := x"2104";
    tmp(64752) := x"2925";
    tmp(64753) := x"2946";
    tmp(64754) := x"3166";
    tmp(64755) := x"3187";
    tmp(64756) := x"3987";
    tmp(64757) := x"39a8";
    tmp(64758) := x"39c8";
    tmp(64759) := x"39c9";
    tmp(64760) := x"39e9";
    tmp(64761) := x"41e9";
    tmp(64762) := x"4209";
    tmp(64763) := x"4209";
    tmp(64764) := x"420a";
    tmp(64765) := x"4a2a";
    tmp(64766) := x"524b";
    tmp(64767) := x"5a6c";
    tmp(64768) := x"5acd";
    tmp(64769) := x"62ce";
    tmp(64770) := x"732f";
    tmp(64771) := x"6b50";
    tmp(64772) := x"7372";
    tmp(64773) := x"83b3";
    tmp(64774) := x"8bf4";
    tmp(64775) := x"8c16";
    tmp(64776) := x"9457";
    tmp(64777) := x"9c98";
    tmp(64778) := x"a4da";
    tmp(64779) := x"ad1b";
    tmp(64780) := x"b57d";
    tmp(64781) := x"bd7d";
    tmp(64782) := x"c5bf";
    tmp(64783) := x"cdff";
    tmp(64784) := x"ce3f";
    tmp(64785) := x"ce3f";
    tmp(64786) := x"ce3f";
    tmp(64787) := x"ce3f";
    tmp(64788) := x"ce3f";
    tmp(64789) := x"c63f";
    tmp(64790) := x"bdfe";
    tmp(64791) := x"b5dd";
    tmp(64792) := x"9d19";
    tmp(64793) := x"94d7";
    tmp(64794) := x"9497";
    tmp(64795) := x"8c76";
    tmp(64796) := x"8414";
    tmp(64797) := x"7bd2";
    tmp(64798) := x"73d2";
    tmp(64799) := x"6bd1";
    tmp(64800) := x"0000";
    tmp(64801) := x"0800";
    tmp(64802) := x"0800";
    tmp(64803) := x"0800";
    tmp(64804) := x"0800";
    tmp(64805) := x"0800";
    tmp(64806) := x"1000";
    tmp(64807) := x"1000";
    tmp(64808) := x"1000";
    tmp(64809) := x"1000";
    tmp(64810) := x"1000";
    tmp(64811) := x"1000";
    tmp(64812) := x"1000";
    tmp(64813) := x"1000";
    tmp(64814) := x"1000";
    tmp(64815) := x"1000";
    tmp(64816) := x"1000";
    tmp(64817) := x"1000";
    tmp(64818) := x"1000";
    tmp(64819) := x"1000";
    tmp(64820) := x"1800";
    tmp(64821) := x"1800";
    tmp(64822) := x"1800";
    tmp(64823) := x"1800";
    tmp(64824) := x"1800";
    tmp(64825) := x"1800";
    tmp(64826) := x"1800";
    tmp(64827) := x"1800";
    tmp(64828) := x"1800";
    tmp(64829) := x"1000";
    tmp(64830) := x"1000";
    tmp(64831) := x"1000";
    tmp(64832) := x"1000";
    tmp(64833) := x"1800";
    tmp(64834) := x"1800";
    tmp(64835) := x"1800";
    tmp(64836) := x"1800";
    tmp(64837) := x"1800";
    tmp(64838) := x"1800";
    tmp(64839) := x"1800";
    tmp(64840) := x"1800";
    tmp(64841) := x"1800";
    tmp(64842) := x"1800";
    tmp(64843) := x"1800";
    tmp(64844) := x"1800";
    tmp(64845) := x"1800";
    tmp(64846) := x"1800";
    tmp(64847) := x"1800";
    tmp(64848) := x"2000";
    tmp(64849) := x"1800";
    tmp(64850) := x"2000";
    tmp(64851) := x"2000";
    tmp(64852) := x"2000";
    tmp(64853) := x"2000";
    tmp(64854) := x"2000";
    tmp(64855) := x"1800";
    tmp(64856) := x"1800";
    tmp(64857) := x"1800";
    tmp(64858) := x"1800";
    tmp(64859) := x"1800";
    tmp(64860) := x"1800";
    tmp(64861) := x"1800";
    tmp(64862) := x"1800";
    tmp(64863) := x"1800";
    tmp(64864) := x"1800";
    tmp(64865) := x"1800";
    tmp(64866) := x"1800";
    tmp(64867) := x"1800";
    tmp(64868) := x"1800";
    tmp(64869) := x"1800";
    tmp(64870) := x"1800";
    tmp(64871) := x"1000";
    tmp(64872) := x"1000";
    tmp(64873) := x"1000";
    tmp(64874) := x"1000";
    tmp(64875) := x"0800";
    tmp(64876) := x"0800";
    tmp(64877) := x"0800";
    tmp(64878) := x"0800";
    tmp(64879) := x"0800";
    tmp(64880) := x"0800";
    tmp(64881) := x"0800";
    tmp(64882) := x"0820";
    tmp(64883) := x"0820";
    tmp(64884) := x"0820";
    tmp(64885) := x"0800";
    tmp(64886) := x"0800";
    tmp(64887) := x"0800";
    tmp(64888) := x"0800";
    tmp(64889) := x"0800";
    tmp(64890) := x"0800";
    tmp(64891) := x"0800";
    tmp(64892) := x"0800";
    tmp(64893) := x"1000";
    tmp(64894) := x"1000";
    tmp(64895) := x"1000";
    tmp(64896) := x"1000";
    tmp(64897) := x"1000";
    tmp(64898) := x"1000";
    tmp(64899) := x"1000";
    tmp(64900) := x"1800";
    tmp(64901) := x"1800";
    tmp(64902) := x"1800";
    tmp(64903) := x"1000";
    tmp(64904) := x"1000";
    tmp(64905) := x"1000";
    tmp(64906) := x"0800";
    tmp(64907) := x"0800";
    tmp(64908) := x"0800";
    tmp(64909) := x"0800";
    tmp(64910) := x"1000";
    tmp(64911) := x"1800";
    tmp(64912) := x"2800";
    tmp(64913) := x"3000";
    tmp(64914) := x"3000";
    tmp(64915) := x"3000";
    tmp(64916) := x"3800";
    tmp(64917) := x"3800";
    tmp(64918) := x"3800";
    tmp(64919) := x"3800";
    tmp(64920) := x"4000";
    tmp(64921) := x"4000";
    tmp(64922) := x"4800";
    tmp(64923) := x"4800";
    tmp(64924) := x"4800";
    tmp(64925) := x"5000";
    tmp(64926) := x"5000";
    tmp(64927) := x"5000";
    tmp(64928) := x"5000";
    tmp(64929) := x"5000";
    tmp(64930) := x"5800";
    tmp(64931) := x"5800";
    tmp(64932) := x"5800";
    tmp(64933) := x"5800";
    tmp(64934) := x"6000";
    tmp(64935) := x"6000";
    tmp(64936) := x"6800";
    tmp(64937) := x"7000";
    tmp(64938) := x"7800";
    tmp(64939) := x"6000";
    tmp(64940) := x"5800";
    tmp(64941) := x"6000";
    tmp(64942) := x"5800";
    tmp(64943) := x"6800";
    tmp(64944) := x"7820";
    tmp(64945) := x"7020";
    tmp(64946) := x"6820";
    tmp(64947) := x"5800";
    tmp(64948) := x"5000";
    tmp(64949) := x"5000";
    tmp(64950) := x"5000";
    tmp(64951) := x"5800";
    tmp(64952) := x"6800";
    tmp(64953) := x"8000";
    tmp(64954) := x"9020";
    tmp(64955) := x"a820";
    tmp(64956) := x"c820";
    tmp(64957) := x"e861";
    tmp(64958) := x"a841";
    tmp(64959) := x"6820";
    tmp(64960) := x"5800";
    tmp(64961) := x"8820";
    tmp(64962) := x"6800";
    tmp(64963) := x"6000";
    tmp(64964) := x"6000";
    tmp(64965) := x"7000";
    tmp(64966) := x"a020";
    tmp(64967) := x"9020";
    tmp(64968) := x"8820";
    tmp(64969) := x"9020";
    tmp(64970) := x"7820";
    tmp(64971) := x"7820";
    tmp(64972) := x"7020";
    tmp(64973) := x"2820";
    tmp(64974) := x"1040";
    tmp(64975) := x"0840";
    tmp(64976) := x"0840";
    tmp(64977) := x"0840";
    tmp(64978) := x"0841";
    tmp(64979) := x"0841";
    tmp(64980) := x"0861";
    tmp(64981) := x"1061";
    tmp(64982) := x"1081";
    tmp(64983) := x"1082";
    tmp(64984) := x"18a2";
    tmp(64985) := x"18c3";
    tmp(64986) := x"18c3";
    tmp(64987) := x"18e4";
    tmp(64988) := x"20e4";
    tmp(64989) := x"2104";
    tmp(64990) := x"2125";
    tmp(64991) := x"2925";
    tmp(64992) := x"2966";
    tmp(64993) := x"3187";
    tmp(64994) := x"3187";
    tmp(64995) := x"39c8";
    tmp(64996) := x"39e9";
    tmp(64997) := x"41e9";
    tmp(64998) := x"420a";
    tmp(64999) := x"4a0a";
    tmp(65000) := x"4a2a";
    tmp(65001) := x"4a4b";
    tmp(65002) := x"4a4b";
    tmp(65003) := x"4a4b";
    tmp(65004) := x"4a4b";
    tmp(65005) := x"526c";
    tmp(65006) := x"5a8d";
    tmp(65007) := x"62ee";
    tmp(65008) := x"6b0f";
    tmp(65009) := x"7351";
    tmp(65010) := x"7b92";
    tmp(65011) := x"7bb2";
    tmp(65012) := x"8bf4";
    tmp(65013) := x"8c15";
    tmp(65014) := x"9457";
    tmp(65015) := x"9cb9";
    tmp(65016) := x"a4da";
    tmp(65017) := x"ad1b";
    tmp(65018) := x"b55d";
    tmp(65019) := x"b57e";
    tmp(65020) := x"c5df";
    tmp(65021) := x"cdff";
    tmp(65022) := x"d63f";
    tmp(65023) := x"ce3f";
    tmp(65024) := x"ce3f";
    tmp(65025) := x"d69f";
    tmp(65026) := x"d69f";
    tmp(65027) := x"ce5f";
    tmp(65028) := x"c63f";
    tmp(65029) := x"c61e";
    tmp(65030) := x"b5bd";
    tmp(65031) := x"ad7b";
    tmp(65032) := x"9cf9";
    tmp(65033) := x"94d7";
    tmp(65034) := x"8c96";
    tmp(65035) := x"8c55";
    tmp(65036) := x"8414";
    tmp(65037) := x"7bd3";
    tmp(65038) := x"73b2";
    tmp(65039) := x"6bd1";
    tmp(65040) := x"0000";
    tmp(65041) := x"0800";
    tmp(65042) := x"0800";
    tmp(65043) := x"0800";
    tmp(65044) := x"0800";
    tmp(65045) := x"1000";
    tmp(65046) := x"1000";
    tmp(65047) := x"1000";
    tmp(65048) := x"1000";
    tmp(65049) := x"1000";
    tmp(65050) := x"1000";
    tmp(65051) := x"1000";
    tmp(65052) := x"1000";
    tmp(65053) := x"1000";
    tmp(65054) := x"1000";
    tmp(65055) := x"0800";
    tmp(65056) := x"1000";
    tmp(65057) := x"1000";
    tmp(65058) := x"1000";
    tmp(65059) := x"1000";
    tmp(65060) := x"1800";
    tmp(65061) := x"1800";
    tmp(65062) := x"1800";
    tmp(65063) := x"1800";
    tmp(65064) := x"1800";
    tmp(65065) := x"1800";
    tmp(65066) := x"1800";
    tmp(65067) := x"1800";
    tmp(65068) := x"1800";
    tmp(65069) := x"1800";
    tmp(65070) := x"1000";
    tmp(65071) := x"1000";
    tmp(65072) := x"1000";
    tmp(65073) := x"1000";
    tmp(65074) := x"1800";
    tmp(65075) := x"1800";
    tmp(65076) := x"1800";
    tmp(65077) := x"1800";
    tmp(65078) := x"1800";
    tmp(65079) := x"1800";
    tmp(65080) := x"1800";
    tmp(65081) := x"1800";
    tmp(65082) := x"1800";
    tmp(65083) := x"1800";
    tmp(65084) := x"1800";
    tmp(65085) := x"1800";
    tmp(65086) := x"1800";
    tmp(65087) := x"1800";
    tmp(65088) := x"1800";
    tmp(65089) := x"1800";
    tmp(65090) := x"1800";
    tmp(65091) := x"1800";
    tmp(65092) := x"2000";
    tmp(65093) := x"1800";
    tmp(65094) := x"1800";
    tmp(65095) := x"1800";
    tmp(65096) := x"1800";
    tmp(65097) := x"1800";
    tmp(65098) := x"1800";
    tmp(65099) := x"1800";
    tmp(65100) := x"1800";
    tmp(65101) := x"1800";
    tmp(65102) := x"1000";
    tmp(65103) := x"1000";
    tmp(65104) := x"1000";
    tmp(65105) := x"1000";
    tmp(65106) := x"1000";
    tmp(65107) := x"1000";
    tmp(65108) := x"1000";
    tmp(65109) := x"1000";
    tmp(65110) := x"1000";
    tmp(65111) := x"1000";
    tmp(65112) := x"1000";
    tmp(65113) := x"1000";
    tmp(65114) := x"0800";
    tmp(65115) := x"0800";
    tmp(65116) := x"0800";
    tmp(65117) := x"0800";
    tmp(65118) := x"0800";
    tmp(65119) := x"0000";
    tmp(65120) := x"0000";
    tmp(65121) := x"0000";
    tmp(65122) := x"0800";
    tmp(65123) := x"0820";
    tmp(65124) := x"0800";
    tmp(65125) := x"0800";
    tmp(65126) := x"0800";
    tmp(65127) := x"0800";
    tmp(65128) := x"0800";
    tmp(65129) := x"0800";
    tmp(65130) := x"0800";
    tmp(65131) := x"0800";
    tmp(65132) := x"0800";
    tmp(65133) := x"0800";
    tmp(65134) := x"1000";
    tmp(65135) := x"1000";
    tmp(65136) := x"1000";
    tmp(65137) := x"1000";
    tmp(65138) := x"1000";
    tmp(65139) := x"1000";
    tmp(65140) := x"1000";
    tmp(65141) := x"1000";
    tmp(65142) := x"1000";
    tmp(65143) := x"1000";
    tmp(65144) := x"1000";
    tmp(65145) := x"1000";
    tmp(65146) := x"0800";
    tmp(65147) := x"0800";
    tmp(65148) := x"0800";
    tmp(65149) := x"1000";
    tmp(65150) := x"1800";
    tmp(65151) := x"2800";
    tmp(65152) := x"3000";
    tmp(65153) := x"3000";
    tmp(65154) := x"3000";
    tmp(65155) := x"3000";
    tmp(65156) := x"3800";
    tmp(65157) := x"3800";
    tmp(65158) := x"3800";
    tmp(65159) := x"3800";
    tmp(65160) := x"3800";
    tmp(65161) := x"4000";
    tmp(65162) := x"4800";
    tmp(65163) := x"4000";
    tmp(65164) := x"5000";
    tmp(65165) := x"5000";
    tmp(65166) := x"5000";
    tmp(65167) := x"5000";
    tmp(65168) := x"5000";
    tmp(65169) := x"5000";
    tmp(65170) := x"5800";
    tmp(65171) := x"5800";
    tmp(65172) := x"5800";
    tmp(65173) := x"6000";
    tmp(65174) := x"6000";
    tmp(65175) := x"6000";
    tmp(65176) := x"7000";
    tmp(65177) := x"7000";
    tmp(65178) := x"7000";
    tmp(65179) := x"6800";
    tmp(65180) := x"6000";
    tmp(65181) := x"5800";
    tmp(65182) := x"5800";
    tmp(65183) := x"6820";
    tmp(65184) := x"6820";
    tmp(65185) := x"6000";
    tmp(65186) := x"6000";
    tmp(65187) := x"5000";
    tmp(65188) := x"5000";
    tmp(65189) := x"4000";
    tmp(65190) := x"4000";
    tmp(65191) := x"6000";
    tmp(65192) := x"7000";
    tmp(65193) := x"8820";
    tmp(65194) := x"a020";
    tmp(65195) := x"b020";
    tmp(65196) := x"c841";
    tmp(65197) := x"d861";
    tmp(65198) := x"9020";
    tmp(65199) := x"6000";
    tmp(65200) := x"5000";
    tmp(65201) := x"7000";
    tmp(65202) := x"6800";
    tmp(65203) := x"5800";
    tmp(65204) := x"5800";
    tmp(65205) := x"8020";
    tmp(65206) := x"9820";
    tmp(65207) := x"8820";
    tmp(65208) := x"9020";
    tmp(65209) := x"9020";
    tmp(65210) := x"7020";
    tmp(65211) := x"6820";
    tmp(65212) := x"4820";
    tmp(65213) := x"1840";
    tmp(65214) := x"0840";
    tmp(65215) := x"0840";
    tmp(65216) := x"0840";
    tmp(65217) := x"0840";
    tmp(65218) := x"0841";
    tmp(65219) := x"0841";
    tmp(65220) := x"0861";
    tmp(65221) := x"1061";
    tmp(65222) := x"1082";
    tmp(65223) := x"10a2";
    tmp(65224) := x"18c2";
    tmp(65225) := x"18c3";
    tmp(65226) := x"18e3";
    tmp(65227) := x"2104";
    tmp(65228) := x"2104";
    tmp(65229) := x"2125";
    tmp(65230) := x"2925";
    tmp(65231) := x"3146";
    tmp(65232) := x"3187";
    tmp(65233) := x"39a8";
    tmp(65234) := x"39e9";
    tmp(65235) := x"41e9";
    tmp(65236) := x"420a";
    tmp(65237) := x"4a2a";
    tmp(65238) := x"4a2b";
    tmp(65239) := x"4a4b";
    tmp(65240) := x"524b";
    tmp(65241) := x"526c";
    tmp(65242) := x"528d";
    tmp(65243) := x"528d";
    tmp(65244) := x"5a8d";
    tmp(65245) := x"62ce";
    tmp(65246) := x"62ef";
    tmp(65247) := x"7331";
    tmp(65248) := x"7b92";
    tmp(65249) := x"7bd4";
    tmp(65250) := x"83d5";
    tmp(65251) := x"8c15";
    tmp(65252) := x"9456";
    tmp(65253) := x"9c77";
    tmp(65254) := x"a4d9";
    tmp(65255) := x"a4fb";
    tmp(65256) := x"b55c";
    tmp(65257) := x"b57d";
    tmp(65258) := x"c5df";
    tmp(65259) := x"c5ff";
    tmp(65260) := x"ce3f";
    tmp(65261) := x"de7f";
    tmp(65262) := x"de9f";
    tmp(65263) := x"de9f";
    tmp(65264) := x"d69f";
    tmp(65265) := x"ce5f";
    tmp(65266) := x"d69f";
    tmp(65267) := x"c63f";
    tmp(65268) := x"c63f";
    tmp(65269) := x"c5fe";
    tmp(65270) := x"b5bc";
    tmp(65271) := x"ad7b";
    tmp(65272) := x"a4f8";
    tmp(65273) := x"9497";
    tmp(65274) := x"9496";
    tmp(65275) := x"8c55";
    tmp(65276) := x"8414";
    tmp(65277) := x"7bd3";
    tmp(65278) := x"7bf3";
    tmp(65279) := x"6bb0";
    tmp(65280) := x"0000";
    tmp(65281) := x"0800";
    tmp(65282) := x"0800";
    tmp(65283) := x"0800";
    tmp(65284) := x"0800";
    tmp(65285) := x"0800";
    tmp(65286) := x"1000";
    tmp(65287) := x"1000";
    tmp(65288) := x"1000";
    tmp(65289) := x"1000";
    tmp(65290) := x"1000";
    tmp(65291) := x"1000";
    tmp(65292) := x"1000";
    tmp(65293) := x"1000";
    tmp(65294) := x"1000";
    tmp(65295) := x"1000";
    tmp(65296) := x"0800";
    tmp(65297) := x"0800";
    tmp(65298) := x"1000";
    tmp(65299) := x"1000";
    tmp(65300) := x"1000";
    tmp(65301) := x"1800";
    tmp(65302) := x"1800";
    tmp(65303) := x"1800";
    tmp(65304) := x"1800";
    tmp(65305) := x"1800";
    tmp(65306) := x"1800";
    tmp(65307) := x"1800";
    tmp(65308) := x"1800";
    tmp(65309) := x"1800";
    tmp(65310) := x"1000";
    tmp(65311) := x"1000";
    tmp(65312) := x"1000";
    tmp(65313) := x"1000";
    tmp(65314) := x"1000";
    tmp(65315) := x"1000";
    tmp(65316) := x"1800";
    tmp(65317) := x"1800";
    tmp(65318) := x"1800";
    tmp(65319) := x"1800";
    tmp(65320) := x"1800";
    tmp(65321) := x"1000";
    tmp(65322) := x"1000";
    tmp(65323) := x"1000";
    tmp(65324) := x"1000";
    tmp(65325) := x"1000";
    tmp(65326) := x"1000";
    tmp(65327) := x"1800";
    tmp(65328) := x"1800";
    tmp(65329) := x"1800";
    tmp(65330) := x"1800";
    tmp(65331) := x"1800";
    tmp(65332) := x"1800";
    tmp(65333) := x"1800";
    tmp(65334) := x"1800";
    tmp(65335) := x"1800";
    tmp(65336) := x"1800";
    tmp(65337) := x"1800";
    tmp(65338) := x"1000";
    tmp(65339) := x"1000";
    tmp(65340) := x"1000";
    tmp(65341) := x"1000";
    tmp(65342) := x"1000";
    tmp(65343) := x"1000";
    tmp(65344) := x"1000";
    tmp(65345) := x"1000";
    tmp(65346) := x"1000";
    tmp(65347) := x"1000";
    tmp(65348) := x"1000";
    tmp(65349) := x"1000";
    tmp(65350) := x"1000";
    tmp(65351) := x"1000";
    tmp(65352) := x"1000";
    tmp(65353) := x"1000";
    tmp(65354) := x"0800";
    tmp(65355) := x"0800";
    tmp(65356) := x"0800";
    tmp(65357) := x"0800";
    tmp(65358) := x"0800";
    tmp(65359) := x"0800";
    tmp(65360) := x"0000";
    tmp(65361) := x"0000";
    tmp(65362) := x"0820";
    tmp(65363) := x"0800";
    tmp(65364) := x"0800";
    tmp(65365) := x"0800";
    tmp(65366) := x"0800";
    tmp(65367) := x"0800";
    tmp(65368) := x"0800";
    tmp(65369) := x"0800";
    tmp(65370) := x"0800";
    tmp(65371) := x"0800";
    tmp(65372) := x"0800";
    tmp(65373) := x"0800";
    tmp(65374) := x"0800";
    tmp(65375) := x"0800";
    tmp(65376) := x"0800";
    tmp(65377) := x"0800";
    tmp(65378) := x"1000";
    tmp(65379) := x"1000";
    tmp(65380) := x"1000";
    tmp(65381) := x"1000";
    tmp(65382) := x"1000";
    tmp(65383) := x"1000";
    tmp(65384) := x"1000";
    tmp(65385) := x"1000";
    tmp(65386) := x"0800";
    tmp(65387) := x"0800";
    tmp(65388) := x"0800";
    tmp(65389) := x"1000";
    tmp(65390) := x"1800";
    tmp(65391) := x"2000";
    tmp(65392) := x"2800";
    tmp(65393) := x"2800";
    tmp(65394) := x"3000";
    tmp(65395) := x"3000";
    tmp(65396) := x"3000";
    tmp(65397) := x"3000";
    tmp(65398) := x"3000";
    tmp(65399) := x"3000";
    tmp(65400) := x"3000";
    tmp(65401) := x"3800";
    tmp(65402) := x"4000";
    tmp(65403) := x"4800";
    tmp(65404) := x"5000";
    tmp(65405) := x"5000";
    tmp(65406) := x"5800";
    tmp(65407) := x"5000";
    tmp(65408) := x"5000";
    tmp(65409) := x"4800";
    tmp(65410) := x"5000";
    tmp(65411) := x"5000";
    tmp(65412) := x"5800";
    tmp(65413) := x"6000";
    tmp(65414) := x"6800";
    tmp(65415) := x"6800";
    tmp(65416) := x"7000";
    tmp(65417) := x"6800";
    tmp(65418) := x"6800";
    tmp(65419) := x"6800";
    tmp(65420) := x"6000";
    tmp(65421) := x"6000";
    tmp(65422) := x"6800";
    tmp(65423) := x"6800";
    tmp(65424) := x"6800";
    tmp(65425) := x"6020";
    tmp(65426) := x"5000";
    tmp(65427) := x"4800";
    tmp(65428) := x"4000";
    tmp(65429) := x"3800";
    tmp(65430) := x"4000";
    tmp(65431) := x"6800";
    tmp(65432) := x"7800";
    tmp(65433) := x"9020";
    tmp(65434) := x"9820";
    tmp(65435) := x"9820";
    tmp(65436) := x"b840";
    tmp(65437) := x"b040";
    tmp(65438) := x"8820";
    tmp(65439) := x"5800";
    tmp(65440) := x"6800";
    tmp(65441) := x"7000";
    tmp(65442) := x"5800";
    tmp(65443) := x"5800";
    tmp(65444) := x"5800";
    tmp(65445) := x"8020";
    tmp(65446) := x"8020";
    tmp(65447) := x"8020";
    tmp(65448) := x"9020";
    tmp(65449) := x"7820";
    tmp(65450) := x"6820";
    tmp(65451) := x"5820";
    tmp(65452) := x"2840";
    tmp(65453) := x"1040";
    tmp(65454) := x"0840";
    tmp(65455) := x"0840";
    tmp(65456) := x"0840";
    tmp(65457) := x"0840";
    tmp(65458) := x"0841";
    tmp(65459) := x"0841";
    tmp(65460) := x"1061";
    tmp(65461) := x"1061";
    tmp(65462) := x"1082";
    tmp(65463) := x"10a2";
    tmp(65464) := x"18c3";
    tmp(65465) := x"18e3";
    tmp(65466) := x"20e4";
    tmp(65467) := x"2104";
    tmp(65468) := x"2125";
    tmp(65469) := x"2925";
    tmp(65470) := x"2946";
    tmp(65471) := x"3186";
    tmp(65472) := x"31a8";
    tmp(65473) := x"39e9";
    tmp(65474) := x"420a";
    tmp(65475) := x"420a";
    tmp(65476) := x"4a2b";
    tmp(65477) := x"4a4b";
    tmp(65478) := x"4a4c";
    tmp(65479) := x"526c";
    tmp(65480) := x"528d";
    tmp(65481) := x"5aad";
    tmp(65482) := x"62ce";
    tmp(65483) := x"62ce";
    tmp(65484) := x"62ef";
    tmp(65485) := x"6b30";
    tmp(65486) := x"7331";
    tmp(65487) := x"7b73";
    tmp(65488) := x"83d5";
    tmp(65489) := x"83f5";
    tmp(65490) := x"8c36";
    tmp(65491) := x"9456";
    tmp(65492) := x"9c77";
    tmp(65493) := x"a4d9";
    tmp(65494) := x"acfa";
    tmp(65495) := x"b55b";
    tmp(65496) := x"bdbe";
    tmp(65497) := x"c5ff";
    tmp(65498) := x"ce3f";
    tmp(65499) := x"d63f";
    tmp(65500) := x"ce3f";
    tmp(65501) := x"d69f";
    tmp(65502) := x"d69f";
    tmp(65503) := x"ce7f";
    tmp(65504) := x"d69f";
    tmp(65505) := x"ce7f";
    tmp(65506) := x"ce7f";
    tmp(65507) := x"c63f";
    tmp(65508) := x"bdfe";
    tmp(65509) := x"b5bc";
    tmp(65510) := x"b5bb";
    tmp(65511) := x"ad79";
    tmp(65512) := x"9cf8";
    tmp(65513) := x"9497";
    tmp(65514) := x"8c55";
    tmp(65515) := x"8434";
    tmp(65516) := x"8434";
    tmp(65517) := x"73b3";
    tmp(65518) := x"73d2";
    tmp(65519) := x"73b1";
    tmp(65520) := x"0000";
    tmp(65521) := x"0800";
    tmp(65522) := x"0800";
    tmp(65523) := x"0800";
    tmp(65524) := x"0800";
    tmp(65525) := x"0800";
    tmp(65526) := x"1000";
    tmp(65527) := x"0800";
    tmp(65528) := x"0800";
    tmp(65529) := x"1000";
    tmp(65530) := x"1000";
    tmp(65531) := x"0800";
    tmp(65532) := x"1000";
    tmp(65533) := x"1000";
    tmp(65534) := x"1000";
    tmp(65535) := x"1000";
    tmp(65536) := x"1000";
    tmp(65537) := x"0800";
    tmp(65538) := x"0800";
    tmp(65539) := x"1000";
    tmp(65540) := x"1000";
    tmp(65541) := x"1800";
    tmp(65542) := x"1800";
    tmp(65543) := x"1800";
    tmp(65544) := x"1800";
    tmp(65545) := x"1800";
    tmp(65546) := x"1800";
    tmp(65547) := x"1800";
    tmp(65548) := x"1800";
    tmp(65549) := x"1800";
    tmp(65550) := x"1800";
    tmp(65551) := x"1000";
    tmp(65552) := x"1000";
    tmp(65553) := x"1000";
    tmp(65554) := x"1000";
    tmp(65555) := x"1000";
    tmp(65556) := x"1000";
    tmp(65557) := x"1000";
    tmp(65558) := x"1000";
    tmp(65559) := x"1000";
    tmp(65560) := x"1000";
    tmp(65561) := x"1000";
    tmp(65562) := x"1000";
    tmp(65563) := x"1000";
    tmp(65564) := x"1000";
    tmp(65565) := x"1000";
    tmp(65566) := x"1000";
    tmp(65567) := x"1000";
    tmp(65568) := x"1800";
    tmp(65569) := x"1800";
    tmp(65570) := x"1800";
    tmp(65571) := x"1800";
    tmp(65572) := x"1800";
    tmp(65573) := x"1800";
    tmp(65574) := x"1800";
    tmp(65575) := x"1800";
    tmp(65576) := x"1000";
    tmp(65577) := x"1000";
    tmp(65578) := x"1000";
    tmp(65579) := x"1000";
    tmp(65580) := x"1000";
    tmp(65581) := x"1000";
    tmp(65582) := x"1000";
    tmp(65583) := x"1000";
    tmp(65584) := x"1000";
    tmp(65585) := x"1000";
    tmp(65586) := x"0800";
    tmp(65587) := x"0800";
    tmp(65588) := x"0800";
    tmp(65589) := x"0800";
    tmp(65590) := x"0800";
    tmp(65591) := x"0800";
    tmp(65592) := x"1000";
    tmp(65593) := x"0800";
    tmp(65594) := x"0800";
    tmp(65595) := x"0800";
    tmp(65596) := x"0800";
    tmp(65597) := x"0800";
    tmp(65598) := x"0800";
    tmp(65599) := x"0000";
    tmp(65600) := x"0000";
    tmp(65601) := x"0000";
    tmp(65602) := x"0800";
    tmp(65603) := x"0800";
    tmp(65604) := x"0800";
    tmp(65605) := x"0800";
    tmp(65606) := x"0800";
    tmp(65607) := x"0800";
    tmp(65608) := x"0800";
    tmp(65609) := x"0800";
    tmp(65610) := x"0800";
    tmp(65611) := x"0800";
    tmp(65612) := x"0800";
    tmp(65613) := x"0800";
    tmp(65614) := x"0800";
    tmp(65615) := x"0800";
    tmp(65616) := x"0800";
    tmp(65617) := x"0800";
    tmp(65618) := x"0800";
    tmp(65619) := x"0800";
    tmp(65620) := x"0800";
    tmp(65621) := x"0800";
    tmp(65622) := x"1000";
    tmp(65623) := x"1000";
    tmp(65624) := x"1000";
    tmp(65625) := x"1000";
    tmp(65626) := x"0800";
    tmp(65627) := x"0800";
    tmp(65628) := x"0800";
    tmp(65629) := x"0800";
    tmp(65630) := x"1000";
    tmp(65631) := x"1000";
    tmp(65632) := x"1800";
    tmp(65633) := x"1800";
    tmp(65634) := x"2000";
    tmp(65635) := x"3000";
    tmp(65636) := x"3000";
    tmp(65637) := x"3000";
    tmp(65638) := x"3000";
    tmp(65639) := x"3000";
    tmp(65640) := x"2800";
    tmp(65641) := x"3000";
    tmp(65642) := x"4000";
    tmp(65643) := x"4800";
    tmp(65644) := x"5000";
    tmp(65645) := x"5800";
    tmp(65646) := x"5800";
    tmp(65647) := x"5000";
    tmp(65648) := x"5000";
    tmp(65649) := x"5000";
    tmp(65650) := x"5000";
    tmp(65651) := x"5000";
    tmp(65652) := x"5800";
    tmp(65653) := x"5800";
    tmp(65654) := x"6000";
    tmp(65655) := x"6800";
    tmp(65656) := x"6800";
    tmp(65657) := x"6800";
    tmp(65658) := x"7020";
    tmp(65659) := x"6800";
    tmp(65660) := x"6000";
    tmp(65661) := x"6000";
    tmp(65662) := x"6800";
    tmp(65663) := x"6800";
    tmp(65664) := x"6820";
    tmp(65665) := x"5820";
    tmp(65666) := x"4800";
    tmp(65667) := x"5000";
    tmp(65668) := x"4000";
    tmp(65669) := x"4000";
    tmp(65670) := x"5000";
    tmp(65671) := x"6800";
    tmp(65672) := x"8020";
    tmp(65673) := x"8820";
    tmp(65674) := x"7800";
    tmp(65675) := x"9020";
    tmp(65676) := x"b020";
    tmp(65677) := x"a020";
    tmp(65678) := x"6800";
    tmp(65679) := x"6800";
    tmp(65680) := x"7820";
    tmp(65681) := x"5800";
    tmp(65682) := x"5800";
    tmp(65683) := x"6000";
    tmp(65684) := x"6000";
    tmp(65685) := x"7820";
    tmp(65686) := x"7820";
    tmp(65687) := x"8020";
    tmp(65688) := x"8020";
    tmp(65689) := x"5820";
    tmp(65690) := x"5040";
    tmp(65691) := x"3840";
    tmp(65692) := x"1040";
    tmp(65693) := x"0840";
    tmp(65694) := x"0840";
    tmp(65695) := x"0840";
    tmp(65696) := x"0840";
    tmp(65697) := x"0840";
    tmp(65698) := x"0841";
    tmp(65699) := x"1061";
    tmp(65700) := x"1061";
    tmp(65701) := x"1081";
    tmp(65702) := x"10a2";
    tmp(65703) := x"18c3";
    tmp(65704) := x"18e3";
    tmp(65705) := x"20e4";
    tmp(65706) := x"2104";
    tmp(65707) := x"2925";
    tmp(65708) := x"2925";
    tmp(65709) := x"2946";
    tmp(65710) := x"3166";
    tmp(65711) := x"3187";
    tmp(65712) := x"39c9";
    tmp(65713) := x"420a";
    tmp(65714) := x"4a2a";
    tmp(65715) := x"4a4b";
    tmp(65716) := x"524c";
    tmp(65717) := x"526d";
    tmp(65718) := x"528d";
    tmp(65719) := x"528d";
    tmp(65720) := x"5aae";
    tmp(65721) := x"62cf";
    tmp(65722) := x"62ef";
    tmp(65723) := x"62ef";
    tmp(65724) := x"6b10";
    tmp(65725) := x"7351";
    tmp(65726) := x"7b93";
    tmp(65727) := x"83d4";
    tmp(65728) := x"8c16";
    tmp(65729) := x"9436";
    tmp(65730) := x"9456";
    tmp(65731) := x"9497";
    tmp(65732) := x"a4d9";
    tmp(65733) := x"ad3b";
    tmp(65734) := x"b55c";
    tmp(65735) := x"bd9d";
    tmp(65736) := x"bdde";
    tmp(65737) := x"c61f";
    tmp(65738) := x"ce3f";
    tmp(65739) := x"d67f";
    tmp(65740) := x"ce7f";
    tmp(65741) := x"d6bf";
    tmp(65742) := x"debf";
    tmp(65743) := x"de9f";
    tmp(65744) := x"ce3f";
    tmp(65745) := x"d65f";
    tmp(65746) := x"d65f";
    tmp(65747) := x"c5ff";
    tmp(65748) := x"bdfe";
    tmp(65749) := x"bddd";
    tmp(65750) := x"b59b";
    tmp(65751) := x"9cf8";
    tmp(65752) := x"9cb7";
    tmp(65753) := x"8c76";
    tmp(65754) := x"8c35";
    tmp(65755) := x"8c54";
    tmp(65756) := x"8414";
    tmp(65757) := x"7bf2";
    tmp(65758) := x"73b1";
    tmp(65759) := x"73b0";
    tmp(65760) := x"0000";
    tmp(65761) := x"0800";
    tmp(65762) := x"0800";
    tmp(65763) := x"0800";
    tmp(65764) := x"0800";
    tmp(65765) := x"0800";
    tmp(65766) := x"0800";
    tmp(65767) := x"0800";
    tmp(65768) := x"0800";
    tmp(65769) := x"0800";
    tmp(65770) := x"0800";
    tmp(65771) := x"0800";
    tmp(65772) := x"1000";
    tmp(65773) := x"1000";
    tmp(65774) := x"1000";
    tmp(65775) := x"1000";
    tmp(65776) := x"1000";
    tmp(65777) := x"0800";
    tmp(65778) := x"1000";
    tmp(65779) := x"1000";
    tmp(65780) := x"1000";
    tmp(65781) := x"1000";
    tmp(65782) := x"1800";
    tmp(65783) := x"1800";
    tmp(65784) := x"1800";
    tmp(65785) := x"1800";
    tmp(65786) := x"1800";
    tmp(65787) := x"1800";
    tmp(65788) := x"1000";
    tmp(65789) := x"1000";
    tmp(65790) := x"1800";
    tmp(65791) := x"1000";
    tmp(65792) := x"1000";
    tmp(65793) := x"1000";
    tmp(65794) := x"1000";
    tmp(65795) := x"1000";
    tmp(65796) := x"0800";
    tmp(65797) := x"1000";
    tmp(65798) := x"1000";
    tmp(65799) := x"1000";
    tmp(65800) := x"1000";
    tmp(65801) := x"1000";
    tmp(65802) := x"1000";
    tmp(65803) := x"1000";
    tmp(65804) := x"1000";
    tmp(65805) := x"1000";
    tmp(65806) := x"1000";
    tmp(65807) := x"1000";
    tmp(65808) := x"1000";
    tmp(65809) := x"1000";
    tmp(65810) := x"1000";
    tmp(65811) := x"1000";
    tmp(65812) := x"1800";
    tmp(65813) := x"1800";
    tmp(65814) := x"1800";
    tmp(65815) := x"1000";
    tmp(65816) := x"1000";
    tmp(65817) := x"1000";
    tmp(65818) := x"1000";
    tmp(65819) := x"1000";
    tmp(65820) := x"1000";
    tmp(65821) := x"1000";
    tmp(65822) := x"0800";
    tmp(65823) := x"0800";
    tmp(65824) := x"0800";
    tmp(65825) := x"0800";
    tmp(65826) := x"0800";
    tmp(65827) := x"0800";
    tmp(65828) := x"0800";
    tmp(65829) := x"0800";
    tmp(65830) := x"0800";
    tmp(65831) := x"0800";
    tmp(65832) := x"1000";
    tmp(65833) := x"0800";
    tmp(65834) := x"0800";
    tmp(65835) := x"0800";
    tmp(65836) := x"0800";
    tmp(65837) := x"0800";
    tmp(65838) := x"0800";
    tmp(65839) := x"0000";
    tmp(65840) := x"0800";
    tmp(65841) := x"0800";
    tmp(65842) := x"0800";
    tmp(65843) := x"0800";
    tmp(65844) := x"0800";
    tmp(65845) := x"0800";
    tmp(65846) := x"0800";
    tmp(65847) := x"0800";
    tmp(65848) := x"0800";
    tmp(65849) := x"0800";
    tmp(65850) := x"0800";
    tmp(65851) := x"0800";
    tmp(65852) := x"0800";
    tmp(65853) := x"0800";
    tmp(65854) := x"0800";
    tmp(65855) := x"0800";
    tmp(65856) := x"0800";
    tmp(65857) := x"0800";
    tmp(65858) := x"0800";
    tmp(65859) := x"0800";
    tmp(65860) := x"0800";
    tmp(65861) := x"0800";
    tmp(65862) := x"0800";
    tmp(65863) := x"0800";
    tmp(65864) := x"0800";
    tmp(65865) := x"0800";
    tmp(65866) := x"0800";
    tmp(65867) := x"0800";
    tmp(65868) := x"0000";
    tmp(65869) := x"0800";
    tmp(65870) := x"0800";
    tmp(65871) := x"0800";
    tmp(65872) := x"0800";
    tmp(65873) := x"1000";
    tmp(65874) := x"2000";
    tmp(65875) := x"3000";
    tmp(65876) := x"3000";
    tmp(65877) := x"3000";
    tmp(65878) := x"3000";
    tmp(65879) := x"3000";
    tmp(65880) := x"3000";
    tmp(65881) := x"2800";
    tmp(65882) := x"4000";
    tmp(65883) := x"5000";
    tmp(65884) := x"5000";
    tmp(65885) := x"5800";
    tmp(65886) := x"5800";
    tmp(65887) := x"5000";
    tmp(65888) := x"5000";
    tmp(65889) := x"5000";
    tmp(65890) := x"5000";
    tmp(65891) := x"5000";
    tmp(65892) := x"5800";
    tmp(65893) := x"5800";
    tmp(65894) := x"6800";
    tmp(65895) := x"6800";
    tmp(65896) := x"6800";
    tmp(65897) := x"6800";
    tmp(65898) := x"7020";
    tmp(65899) := x"6800";
    tmp(65900) := x"6000";
    tmp(65901) := x"6000";
    tmp(65902) := x"6800";
    tmp(65903) := x"7020";
    tmp(65904) := x"6820";
    tmp(65905) := x"5820";
    tmp(65906) := x"5820";
    tmp(65907) := x"4800";
    tmp(65908) := x"4000";
    tmp(65909) := x"5000";
    tmp(65910) := x"6000";
    tmp(65911) := x"7800";
    tmp(65912) := x"7820";
    tmp(65913) := x"6800";
    tmp(65914) := x"7000";
    tmp(65915) := x"9020";
    tmp(65916) := x"a820";
    tmp(65917) := x"8020";
    tmp(65918) := x"6800";
    tmp(65919) := x"8020";
    tmp(65920) := x"6800";
    tmp(65921) := x"5800";
    tmp(65922) := x"7000";
    tmp(65923) := x"6800";
    tmp(65924) := x"7020";
    tmp(65925) := x"8020";
    tmp(65926) := x"7820";
    tmp(65927) := x"7820";
    tmp(65928) := x"5820";
    tmp(65929) := x"2840";
    tmp(65930) := x"2040";
    tmp(65931) := x"1840";
    tmp(65932) := x"0840";
    tmp(65933) := x"0840";
    tmp(65934) := x"0840";
    tmp(65935) := x"0840";
    tmp(65936) := x"0840";
    tmp(65937) := x"0840";
    tmp(65938) := x"1061";
    tmp(65939) := x"1061";
    tmp(65940) := x"1081";
    tmp(65941) := x"10a2";
    tmp(65942) := x"18a2";
    tmp(65943) := x"18c3";
    tmp(65944) := x"20e4";
    tmp(65945) := x"2105";
    tmp(65946) := x"2925";
    tmp(65947) := x"2946";
    tmp(65948) := x"2946";
    tmp(65949) := x"3166";
    tmp(65950) := x"3187";
    tmp(65951) := x"39a8";
    tmp(65952) := x"41ea";
    tmp(65953) := x"420a";
    tmp(65954) := x"4a4b";
    tmp(65955) := x"526c";
    tmp(65956) := x"526d";
    tmp(65957) := x"528d";
    tmp(65958) := x"5a8d";
    tmp(65959) := x"5aae";
    tmp(65960) := x"5acf";
    tmp(65961) := x"62ef";
    tmp(65962) := x"6b30";
    tmp(65963) := x"6b31";
    tmp(65964) := x"6b51";
    tmp(65965) := x"7372";
    tmp(65966) := x"7b93";
    tmp(65967) := x"7bb4";
    tmp(65968) := x"8c16";
    tmp(65969) := x"9477";
    tmp(65970) := x"9477";
    tmp(65971) := x"9c98";
    tmp(65972) := x"acf9";
    tmp(65973) := x"ad3b";
    tmp(65974) := x"b57c";
    tmp(65975) := x"bdbd";
    tmp(65976) := x"c5fe";
    tmp(65977) := x"ce1f";
    tmp(65978) := x"ce1f";
    tmp(65979) := x"ce3f";
    tmp(65980) := x"ce7f";
    tmp(65981) := x"de9f";
    tmp(65982) := x"de9f";
    tmp(65983) := x"d67f";
    tmp(65984) := x"ce5f";
    tmp(65985) := x"d63f";
    tmp(65986) := x"c63f";
    tmp(65987) := x"c5fe";
    tmp(65988) := x"bdbd";
    tmp(65989) := x"b5bd";
    tmp(65990) := x"ad7a";
    tmp(65991) := x"9cd8";
    tmp(65992) := x"9c97";
    tmp(65993) := x"8c55";
    tmp(65994) := x"8c15";
    tmp(65995) := x"8414";
    tmp(65996) := x"8413";
    tmp(65997) := x"7bd2";
    tmp(65998) := x"73b1";
    tmp(65999) := x"6b4f";
    tmp(66000) := x"0000";
    tmp(66001) := x"0800";
    tmp(66002) := x"0800";
    tmp(66003) := x"0800";
    tmp(66004) := x"0800";
    tmp(66005) := x"0800";
    tmp(66006) := x"0800";
    tmp(66007) := x"0800";
    tmp(66008) := x"0800";
    tmp(66009) := x"0800";
    tmp(66010) := x"0800";
    tmp(66011) := x"0800";
    tmp(66012) := x"0800";
    tmp(66013) := x"0800";
    tmp(66014) := x"1000";
    tmp(66015) := x"1000";
    tmp(66016) := x"1000";
    tmp(66017) := x"1000";
    tmp(66018) := x"1000";
    tmp(66019) := x"1000";
    tmp(66020) := x"1000";
    tmp(66021) := x"1000";
    tmp(66022) := x"1000";
    tmp(66023) := x"1000";
    tmp(66024) := x"1000";
    tmp(66025) := x"1000";
    tmp(66026) := x"1800";
    tmp(66027) := x"1800";
    tmp(66028) := x"1000";
    tmp(66029) := x"1000";
    tmp(66030) := x"1000";
    tmp(66031) := x"1000";
    tmp(66032) := x"1000";
    tmp(66033) := x"1000";
    tmp(66034) := x"0800";
    tmp(66035) := x"0800";
    tmp(66036) := x"0800";
    tmp(66037) := x"0800";
    tmp(66038) := x"1000";
    tmp(66039) := x"1000";
    tmp(66040) := x"1000";
    tmp(66041) := x"1000";
    tmp(66042) := x"1000";
    tmp(66043) := x"1000";
    tmp(66044) := x"1000";
    tmp(66045) := x"1000";
    tmp(66046) := x"1000";
    tmp(66047) := x"1000";
    tmp(66048) := x"1000";
    tmp(66049) := x"1000";
    tmp(66050) := x"1000";
    tmp(66051) := x"1000";
    tmp(66052) := x"1000";
    tmp(66053) := x"1000";
    tmp(66054) := x"1000";
    tmp(66055) := x"1000";
    tmp(66056) := x"1000";
    tmp(66057) := x"1000";
    tmp(66058) := x"1000";
    tmp(66059) := x"1000";
    tmp(66060) := x"0800";
    tmp(66061) := x"0800";
    tmp(66062) := x"0800";
    tmp(66063) := x"0800";
    tmp(66064) := x"0800";
    tmp(66065) := x"0800";
    tmp(66066) := x"0800";
    tmp(66067) := x"0800";
    tmp(66068) := x"0800";
    tmp(66069) := x"0800";
    tmp(66070) := x"1000";
    tmp(66071) := x"1000";
    tmp(66072) := x"1000";
    tmp(66073) := x"1000";
    tmp(66074) := x"1000";
    tmp(66075) := x"1000";
    tmp(66076) := x"1820";
    tmp(66077) := x"1820";
    tmp(66078) := x"1821";
    tmp(66079) := x"1821";
    tmp(66080) := x"1020";
    tmp(66081) := x"1020";
    tmp(66082) := x"1000";
    tmp(66083) := x"1000";
    tmp(66084) := x"1000";
    tmp(66085) := x"1000";
    tmp(66086) := x"1800";
    tmp(66087) := x"1820";
    tmp(66088) := x"1000";
    tmp(66089) := x"1000";
    tmp(66090) := x"1000";
    tmp(66091) := x"1800";
    tmp(66092) := x"1000";
    tmp(66093) := x"1000";
    tmp(66094) := x"1020";
    tmp(66095) := x"1020";
    tmp(66096) := x"1000";
    tmp(66097) := x"1000";
    tmp(66098) := x"1000";
    tmp(66099) := x"0800";
    tmp(66100) := x"0800";
    tmp(66101) := x"0800";
    tmp(66102) := x"0800";
    tmp(66103) := x"0800";
    tmp(66104) := x"0000";
    tmp(66105) := x"0000";
    tmp(66106) := x"0000";
    tmp(66107) := x"0000";
    tmp(66108) := x"0000";
    tmp(66109) := x"0000";
    tmp(66110) := x"0000";
    tmp(66111) := x"0000";
    tmp(66112) := x"0800";
    tmp(66113) := x"1000";
    tmp(66114) := x"2000";
    tmp(66115) := x"2800";
    tmp(66116) := x"2800";
    tmp(66117) := x"3000";
    tmp(66118) := x"3000";
    tmp(66119) := x"2800";
    tmp(66120) := x"3000";
    tmp(66121) := x"3800";
    tmp(66122) := x"4800";
    tmp(66123) := x"5000";
    tmp(66124) := x"5800";
    tmp(66125) := x"5800";
    tmp(66126) := x"5800";
    tmp(66127) := x"5000";
    tmp(66128) := x"5000";
    tmp(66129) := x"4800";
    tmp(66130) := x"5000";
    tmp(66131) := x"5800";
    tmp(66132) := x"5800";
    tmp(66133) := x"6000";
    tmp(66134) := x"6820";
    tmp(66135) := x"6800";
    tmp(66136) := x"6000";
    tmp(66137) := x"6800";
    tmp(66138) := x"7000";
    tmp(66139) := x"6800";
    tmp(66140) := x"6800";
    tmp(66141) := x"6000";
    tmp(66142) := x"6820";
    tmp(66143) := x"7020";
    tmp(66144) := x"6820";
    tmp(66145) := x"7020";
    tmp(66146) := x"6820";
    tmp(66147) := x"5000";
    tmp(66148) := x"5000";
    tmp(66149) := x"5800";
    tmp(66150) := x"7000";
    tmp(66151) := x"7800";
    tmp(66152) := x"6000";
    tmp(66153) := x"5800";
    tmp(66154) := x"7800";
    tmp(66155) := x"8820";
    tmp(66156) := x"9020";
    tmp(66157) := x"6800";
    tmp(66158) := x"7000";
    tmp(66159) := x"7000";
    tmp(66160) := x"5800";
    tmp(66161) := x"7800";
    tmp(66162) := x"8820";
    tmp(66163) := x"7000";
    tmp(66164) := x"7820";
    tmp(66165) := x"7820";
    tmp(66166) := x"7820";
    tmp(66167) := x"5820";
    tmp(66168) := x"2840";
    tmp(66169) := x"1041";
    tmp(66170) := x"1041";
    tmp(66171) := x"0840";
    tmp(66172) := x"0840";
    tmp(66173) := x"0840";
    tmp(66174) := x"0840";
    tmp(66175) := x"0840";
    tmp(66176) := x"0840";
    tmp(66177) := x"0841";
    tmp(66178) := x"1061";
    tmp(66179) := x"1061";
    tmp(66180) := x"1081";
    tmp(66181) := x"10a2";
    tmp(66182) := x"18a2";
    tmp(66183) := x"18e3";
    tmp(66184) := x"2104";
    tmp(66185) := x"2925";
    tmp(66186) := x"2946";
    tmp(66187) := x"2946";
    tmp(66188) := x"3167";
    tmp(66189) := x"3187";
    tmp(66190) := x"39c8";
    tmp(66191) := x"39c9";
    tmp(66192) := x"420a";
    tmp(66193) := x"422b";
    tmp(66194) := x"4a4c";
    tmp(66195) := x"4a4c";
    tmp(66196) := x"528d";
    tmp(66197) := x"528d";
    tmp(66198) := x"528e";
    tmp(66199) := x"5ace";
    tmp(66200) := x"62cf";
    tmp(66201) := x"62f0";
    tmp(66202) := x"6b11";
    tmp(66203) := x"6b30";
    tmp(66204) := x"7352";
    tmp(66205) := x"7393";
    tmp(66206) := x"7bb4";
    tmp(66207) := x"83f5";
    tmp(66208) := x"8c16";
    tmp(66209) := x"9477";
    tmp(66210) := x"9c77";
    tmp(66211) := x"a4b9";
    tmp(66212) := x"acfa";
    tmp(66213) := x"b55c";
    tmp(66214) := x"bd9d";
    tmp(66215) := x"c5be";
    tmp(66216) := x"c5ff";
    tmp(66217) := x"ce3f";
    tmp(66218) := x"ce3f";
    tmp(66219) := x"ce5f";
    tmp(66220) := x"d67f";
    tmp(66221) := x"de7f";
    tmp(66222) := x"de9f";
    tmp(66223) := x"d67f";
    tmp(66224) := x"c61f";
    tmp(66225) := x"ce3f";
    tmp(66226) := x"bdfe";
    tmp(66227) := x"bdbd";
    tmp(66228) := x"b57c";
    tmp(66229) := x"b57b";
    tmp(66230) := x"a519";
    tmp(66231) := x"94d7";
    tmp(66232) := x"9496";
    tmp(66233) := x"8c56";
    tmp(66234) := x"8c15";
    tmp(66235) := x"83f4";
    tmp(66236) := x"8413";
    tmp(66237) := x"7bd2";
    tmp(66238) := x"7390";
    tmp(66239) := x"6b4f";
    tmp(66240) := x"0000";
    tmp(66241) := x"0800";
    tmp(66242) := x"0800";
    tmp(66243) := x"0800";
    tmp(66244) := x"0800";
    tmp(66245) := x"0800";
    tmp(66246) := x"0800";
    tmp(66247) := x"0800";
    tmp(66248) := x"0800";
    tmp(66249) := x"0800";
    tmp(66250) := x"0800";
    tmp(66251) := x"0800";
    tmp(66252) := x"0800";
    tmp(66253) := x"0800";
    tmp(66254) := x"0800";
    tmp(66255) := x"0800";
    tmp(66256) := x"0800";
    tmp(66257) := x"1000";
    tmp(66258) := x"1000";
    tmp(66259) := x"1000";
    tmp(66260) := x"1000";
    tmp(66261) := x"1000";
    tmp(66262) := x"1000";
    tmp(66263) := x"1000";
    tmp(66264) := x"1000";
    tmp(66265) := x"1000";
    tmp(66266) := x"1000";
    tmp(66267) := x"1000";
    tmp(66268) := x"1000";
    tmp(66269) := x"1000";
    tmp(66270) := x"1000";
    tmp(66271) := x"1000";
    tmp(66272) := x"1000";
    tmp(66273) := x"0800";
    tmp(66274) := x"0800";
    tmp(66275) := x"0800";
    tmp(66276) := x"0800";
    tmp(66277) := x"0800";
    tmp(66278) := x"0800";
    tmp(66279) := x"0800";
    tmp(66280) := x"0800";
    tmp(66281) := x"0800";
    tmp(66282) := x"1000";
    tmp(66283) := x"1000";
    tmp(66284) := x"1000";
    tmp(66285) := x"1000";
    tmp(66286) := x"1000";
    tmp(66287) := x"1000";
    tmp(66288) := x"1000";
    tmp(66289) := x"1000";
    tmp(66290) := x"1000";
    tmp(66291) := x"1000";
    tmp(66292) := x"1000";
    tmp(66293) := x"0800";
    tmp(66294) := x"0800";
    tmp(66295) := x"0800";
    tmp(66296) := x"0800";
    tmp(66297) := x"0800";
    tmp(66298) := x"0800";
    tmp(66299) := x"0800";
    tmp(66300) := x"0800";
    tmp(66301) := x"0800";
    tmp(66302) := x"1000";
    tmp(66303) := x"1000";
    tmp(66304) := x"1800";
    tmp(66305) := x"2020";
    tmp(66306) := x"2820";
    tmp(66307) := x"3041";
    tmp(66308) := x"3041";
    tmp(66309) := x"2020";
    tmp(66310) := x"1000";
    tmp(66311) := x"1000";
    tmp(66312) := x"1020";
    tmp(66313) := x"1020";
    tmp(66314) := x"1020";
    tmp(66315) := x"0820";
    tmp(66316) := x"1020";
    tmp(66317) := x"1021";
    tmp(66318) := x"1841";
    tmp(66319) := x"1841";
    tmp(66320) := x"1820";
    tmp(66321) := x"1020";
    tmp(66322) := x"0800";
    tmp(66323) := x"0820";
    tmp(66324) := x"0820";
    tmp(66325) := x"1020";
    tmp(66326) := x"1020";
    tmp(66327) := x"1820";
    tmp(66328) := x"1020";
    tmp(66329) := x"0820";
    tmp(66330) := x"1020";
    tmp(66331) := x"1000";
    tmp(66332) := x"0800";
    tmp(66333) := x"0800";
    tmp(66334) := x"0800";
    tmp(66335) := x"0800";
    tmp(66336) := x"1000";
    tmp(66337) := x"1800";
    tmp(66338) := x"1000";
    tmp(66339) := x"1000";
    tmp(66340) := x"1020";
    tmp(66341) := x"1000";
    tmp(66342) := x"1000";
    tmp(66343) := x"1000";
    tmp(66344) := x"0800";
    tmp(66345) := x"0800";
    tmp(66346) := x"0000";
    tmp(66347) := x"0000";
    tmp(66348) := x"0000";
    tmp(66349) := x"0800";
    tmp(66350) := x"0800";
    tmp(66351) := x"0800";
    tmp(66352) := x"1000";
    tmp(66353) := x"1000";
    tmp(66354) := x"1800";
    tmp(66355) := x"2800";
    tmp(66356) := x"2800";
    tmp(66357) := x"2800";
    tmp(66358) := x"3000";
    tmp(66359) := x"3000";
    tmp(66360) := x"3800";
    tmp(66361) := x"4800";
    tmp(66362) := x"4800";
    tmp(66363) := x"5000";
    tmp(66364) := x"5000";
    tmp(66365) := x"6000";
    tmp(66366) := x"5000";
    tmp(66367) := x"4000";
    tmp(66368) := x"4800";
    tmp(66369) := x"4800";
    tmp(66370) := x"5000";
    tmp(66371) := x"5800";
    tmp(66372) := x"5800";
    tmp(66373) := x"6000";
    tmp(66374) := x"6000";
    tmp(66375) := x"6000";
    tmp(66376) := x"5800";
    tmp(66377) := x"6800";
    tmp(66378) := x"6800";
    tmp(66379) := x"6800";
    tmp(66380) := x"6800";
    tmp(66381) := x"6000";
    tmp(66382) := x"7020";
    tmp(66383) := x"7820";
    tmp(66384) := x"7820";
    tmp(66385) := x"7821";
    tmp(66386) := x"6820";
    tmp(66387) := x"5820";
    tmp(66388) := x"5000";
    tmp(66389) := x"6000";
    tmp(66390) := x"6800";
    tmp(66391) := x"6800";
    tmp(66392) := x"5000";
    tmp(66393) := x"7000";
    tmp(66394) := x"7800";
    tmp(66395) := x"8820";
    tmp(66396) := x"7000";
    tmp(66397) := x"7000";
    tmp(66398) := x"7000";
    tmp(66399) := x"5800";
    tmp(66400) := x"7000";
    tmp(66401) := x"8820";
    tmp(66402) := x"8820";
    tmp(66403) := x"6800";
    tmp(66404) := x"7020";
    tmp(66405) := x"6820";
    tmp(66406) := x"5820";
    tmp(66407) := x"2840";
    tmp(66408) := x"1061";
    tmp(66409) := x"1061";
    tmp(66410) := x"1061";
    tmp(66411) := x"0841";
    tmp(66412) := x"0840";
    tmp(66413) := x"0840";
    tmp(66414) := x"0840";
    tmp(66415) := x"0840";
    tmp(66416) := x"0840";
    tmp(66417) := x"0840";
    tmp(66418) := x"0841";
    tmp(66419) := x"1061";
    tmp(66420) := x"1081";
    tmp(66421) := x"10a2";
    tmp(66422) := x"18a2";
    tmp(66423) := x"18e3";
    tmp(66424) := x"2104";
    tmp(66425) := x"2125";
    tmp(66426) := x"2946";
    tmp(66427) := x"2966";
    tmp(66428) := x"3187";
    tmp(66429) := x"31a8";
    tmp(66430) := x"39c9";
    tmp(66431) := x"39ea";
    tmp(66432) := x"422a";
    tmp(66433) := x"4a2b";
    tmp(66434) := x"524c";
    tmp(66435) := x"526c";
    tmp(66436) := x"526c";
    tmp(66437) := x"528d";
    tmp(66438) := x"5a8e";
    tmp(66439) := x"5aae";
    tmp(66440) := x"5acf";
    tmp(66441) := x"62f0";
    tmp(66442) := x"6310";
    tmp(66443) := x"6b51";
    tmp(66444) := x"7372";
    tmp(66445) := x"7372";
    tmp(66446) := x"7bb4";
    tmp(66447) := x"83f5";
    tmp(66448) := x"9477";
    tmp(66449) := x"9478";
    tmp(66450) := x"9cb9";
    tmp(66451) := x"9c99";
    tmp(66452) := x"ad3b";
    tmp(66453) := x"b55d";
    tmp(66454) := x"bd9e";
    tmp(66455) := x"c5df";
    tmp(66456) := x"cdff";
    tmp(66457) := x"ce3f";
    tmp(66458) := x"ce5f";
    tmp(66459) := x"d69f";
    tmp(66460) := x"de9f";
    tmp(66461) := x"de9f";
    tmp(66462) := x"ce5f";
    tmp(66463) := x"ce5f";
    tmp(66464) := x"ce3f";
    tmp(66465) := x"be1e";
    tmp(66466) := x"bdfd";
    tmp(66467) := x"bd9d";
    tmp(66468) := x"b53b";
    tmp(66469) := x"ad3a";
    tmp(66470) := x"9cd8";
    tmp(66471) := x"8c76";
    tmp(66472) := x"8c55";
    tmp(66473) := x"8454";
    tmp(66474) := x"8c14";
    tmp(66475) := x"7bd3";
    tmp(66476) := x"7bf3";
    tmp(66477) := x"73b0";
    tmp(66478) := x"6b6e";
    tmp(66479) := x"6b4e";
    tmp(66480) := x"0000";
    tmp(66481) := x"0800";
    tmp(66482) := x"0800";
    tmp(66483) := x"0800";
    tmp(66484) := x"0800";
    tmp(66485) := x"0800";
    tmp(66486) := x"0800";
    tmp(66487) := x"0800";
    tmp(66488) := x"0800";
    tmp(66489) := x"0800";
    tmp(66490) := x"0800";
    tmp(66491) := x"0800";
    tmp(66492) := x"0800";
    tmp(66493) := x"0800";
    tmp(66494) := x"1000";
    tmp(66495) := x"1000";
    tmp(66496) := x"1000";
    tmp(66497) := x"1000";
    tmp(66498) := x"1000";
    tmp(66499) := x"1000";
    tmp(66500) := x"1000";
    tmp(66501) := x"1000";
    tmp(66502) := x"1000";
    tmp(66503) := x"1000";
    tmp(66504) := x"1000";
    tmp(66505) := x"1000";
    tmp(66506) := x"1000";
    tmp(66507) := x"1000";
    tmp(66508) := x"1000";
    tmp(66509) := x"1000";
    tmp(66510) := x"1000";
    tmp(66511) := x"0800";
    tmp(66512) := x"0800";
    tmp(66513) := x"0800";
    tmp(66514) := x"0800";
    tmp(66515) := x"0800";
    tmp(66516) := x"0800";
    tmp(66517) := x"0800";
    tmp(66518) := x"0800";
    tmp(66519) := x"0800";
    tmp(66520) := x"1000";
    tmp(66521) := x"1000";
    tmp(66522) := x"1000";
    tmp(66523) := x"1000";
    tmp(66524) := x"1000";
    tmp(66525) := x"1000";
    tmp(66526) := x"1000";
    tmp(66527) := x"0800";
    tmp(66528) := x"1000";
    tmp(66529) := x"0800";
    tmp(66530) := x"0800";
    tmp(66531) := x"0800";
    tmp(66532) := x"0800";
    tmp(66533) := x"0800";
    tmp(66534) := x"1000";
    tmp(66535) := x"1000";
    tmp(66536) := x"1000";
    tmp(66537) := x"1800";
    tmp(66538) := x"1800";
    tmp(66539) := x"2020";
    tmp(66540) := x"2820";
    tmp(66541) := x"2820";
    tmp(66542) := x"2820";
    tmp(66543) := x"2841";
    tmp(66544) := x"2841";
    tmp(66545) := x"2841";
    tmp(66546) := x"2841";
    tmp(66547) := x"2820";
    tmp(66548) := x"2020";
    tmp(66549) := x"2020";
    tmp(66550) := x"1820";
    tmp(66551) := x"1841";
    tmp(66552) := x"1041";
    tmp(66553) := x"0840";
    tmp(66554) := x"0820";
    tmp(66555) := x"0820";
    tmp(66556) := x"0820";
    tmp(66557) := x"0820";
    tmp(66558) := x"0840";
    tmp(66559) := x"0820";
    tmp(66560) := x"0820";
    tmp(66561) := x"0800";
    tmp(66562) := x"0800";
    tmp(66563) := x"0820";
    tmp(66564) := x"0820";
    tmp(66565) := x"0820";
    tmp(66566) := x"0841";
    tmp(66567) := x"0841";
    tmp(66568) := x"0841";
    tmp(66569) := x"0841";
    tmp(66570) := x"0841";
    tmp(66571) := x"0820";
    tmp(66572) := x"0800";
    tmp(66573) := x"0800";
    tmp(66574) := x"0800";
    tmp(66575) := x"0800";
    tmp(66576) := x"1000";
    tmp(66577) := x"1820";
    tmp(66578) := x"2020";
    tmp(66579) := x"1820";
    tmp(66580) := x"1020";
    tmp(66581) := x"1020";
    tmp(66582) := x"1020";
    tmp(66583) := x"1800";
    tmp(66584) := x"1000";
    tmp(66585) := x"0800";
    tmp(66586) := x"0800";
    tmp(66587) := x"0800";
    tmp(66588) := x"0000";
    tmp(66589) := x"0000";
    tmp(66590) := x"0800";
    tmp(66591) := x"0800";
    tmp(66592) := x"1000";
    tmp(66593) := x"1000";
    tmp(66594) := x"1800";
    tmp(66595) := x"2000";
    tmp(66596) := x"2800";
    tmp(66597) := x"2800";
    tmp(66598) := x"3000";
    tmp(66599) := x"3000";
    tmp(66600) := x"3800";
    tmp(66601) := x"4800";
    tmp(66602) := x"5000";
    tmp(66603) := x"5000";
    tmp(66604) := x"5800";
    tmp(66605) := x"6000";
    tmp(66606) := x"5000";
    tmp(66607) := x"4800";
    tmp(66608) := x"3800";
    tmp(66609) := x"3000";
    tmp(66610) := x"4000";
    tmp(66611) := x"5000";
    tmp(66612) := x"5000";
    tmp(66613) := x"5800";
    tmp(66614) := x"5800";
    tmp(66615) := x"5800";
    tmp(66616) := x"6800";
    tmp(66617) := x"6800";
    tmp(66618) := x"6800";
    tmp(66619) := x"6800";
    tmp(66620) := x"5800";
    tmp(66621) := x"6820";
    tmp(66622) := x"8020";
    tmp(66623) := x"7020";
    tmp(66624) := x"7820";
    tmp(66625) := x"7820";
    tmp(66626) := x"6820";
    tmp(66627) := x"5000";
    tmp(66628) := x"5800";
    tmp(66629) := x"6000";
    tmp(66630) := x"6000";
    tmp(66631) := x"5000";
    tmp(66632) := x"6000";
    tmp(66633) := x"6800";
    tmp(66634) := x"7800";
    tmp(66635) := x"7800";
    tmp(66636) := x"7000";
    tmp(66637) := x"7000";
    tmp(66638) := x"6000";
    tmp(66639) := x"6000";
    tmp(66640) := x"8020";
    tmp(66641) := x"8820";
    tmp(66642) := x"6800";
    tmp(66643) := x"6000";
    tmp(66644) := x"6020";
    tmp(66645) := x"5840";
    tmp(66646) := x"3040";
    tmp(66647) := x"1861";
    tmp(66648) := x"1061";
    tmp(66649) := x"1061";
    tmp(66650) := x"1061";
    tmp(66651) := x"1061";
    tmp(66652) := x"0841";
    tmp(66653) := x"0840";
    tmp(66654) := x"0840";
    tmp(66655) := x"0840";
    tmp(66656) := x"0840";
    tmp(66657) := x"0840";
    tmp(66658) := x"0840";
    tmp(66659) := x"1061";
    tmp(66660) := x"1061";
    tmp(66661) := x"10a2";
    tmp(66662) := x"18a2";
    tmp(66663) := x"18c3";
    tmp(66664) := x"20e4";
    tmp(66665) := x"2104";
    tmp(66666) := x"2925";
    tmp(66667) := x"2946";
    tmp(66668) := x"3187";
    tmp(66669) := x"31a8";
    tmp(66670) := x"39c9";
    tmp(66671) := x"39ea";
    tmp(66672) := x"420a";
    tmp(66673) := x"4a4b";
    tmp(66674) := x"4a4b";
    tmp(66675) := x"4a4c";
    tmp(66676) := x"526d";
    tmp(66677) := x"528d";
    tmp(66678) := x"528d";
    tmp(66679) := x"5aae";
    tmp(66680) := x"62ef";
    tmp(66681) := x"62ef";
    tmp(66682) := x"6310";
    tmp(66683) := x"6b31";
    tmp(66684) := x"7372";
    tmp(66685) := x"7b93";
    tmp(66686) := x"7bd4";
    tmp(66687) := x"83f5";
    tmp(66688) := x"9457";
    tmp(66689) := x"9479";
    tmp(66690) := x"9499";
    tmp(66691) := x"a4fa";
    tmp(66692) := x"b55c";
    tmp(66693) := x"bd9d";
    tmp(66694) := x"c5df";
    tmp(66695) := x"ce3f";
    tmp(66696) := x"d63f";
    tmp(66697) := x"ce3f";
    tmp(66698) := x"ce3f";
    tmp(66699) := x"ce3f";
    tmp(66700) := x"ce5f";
    tmp(66701) := x"de9f";
    tmp(66702) := x"d67f";
    tmp(66703) := x"ce3f";
    tmp(66704) := x"c5de";
    tmp(66705) := x"bdbe";
    tmp(66706) := x"bdbd";
    tmp(66707) := x"b55b";
    tmp(66708) := x"ad3a";
    tmp(66709) := x"a4f9";
    tmp(66710) := x"94d8";
    tmp(66711) := x"9496";
    tmp(66712) := x"8c55";
    tmp(66713) := x"8413";
    tmp(66714) := x"83d2";
    tmp(66715) := x"7bd2";
    tmp(66716) := x"7bb1";
    tmp(66717) := x"6b90";
    tmp(66718) := x"6b4e";
    tmp(66719) := x"632e";
    tmp(66720) := x"0000";
    tmp(66721) := x"0800";
    tmp(66722) := x"0800";
    tmp(66723) := x"0800";
    tmp(66724) := x"0800";
    tmp(66725) := x"0800";
    tmp(66726) := x"0800";
    tmp(66727) := x"0800";
    tmp(66728) := x"0800";
    tmp(66729) := x"0800";
    tmp(66730) := x"0800";
    tmp(66731) := x"0800";
    tmp(66732) := x"0800";
    tmp(66733) := x"0800";
    tmp(66734) := x"0800";
    tmp(66735) := x"0800";
    tmp(66736) := x"0800";
    tmp(66737) := x"1000";
    tmp(66738) := x"1000";
    tmp(66739) := x"1000";
    tmp(66740) := x"1000";
    tmp(66741) := x"1000";
    tmp(66742) := x"1000";
    tmp(66743) := x"0800";
    tmp(66744) := x"1000";
    tmp(66745) := x"1000";
    tmp(66746) := x"1000";
    tmp(66747) := x"1000";
    tmp(66748) := x"0800";
    tmp(66749) := x"0800";
    tmp(66750) := x"0800";
    tmp(66751) := x"0800";
    tmp(66752) := x"0800";
    tmp(66753) := x"0800";
    tmp(66754) := x"0800";
    tmp(66755) := x"1000";
    tmp(66756) := x"1000";
    tmp(66757) := x"1000";
    tmp(66758) := x"1000";
    tmp(66759) := x"1000";
    tmp(66760) := x"1000";
    tmp(66761) := x"1000";
    tmp(66762) := x"1000";
    tmp(66763) := x"1000";
    tmp(66764) := x"1000";
    tmp(66765) := x"1000";
    tmp(66766) := x"1000";
    tmp(66767) := x"1000";
    tmp(66768) := x"1000";
    tmp(66769) := x"1000";
    tmp(66770) := x"1000";
    tmp(66771) := x"1000";
    tmp(66772) := x"1800";
    tmp(66773) := x"2000";
    tmp(66774) := x"2820";
    tmp(66775) := x"2820";
    tmp(66776) := x"2820";
    tmp(66777) := x"2820";
    tmp(66778) := x"3041";
    tmp(66779) := x"2821";
    tmp(66780) := x"2021";
    tmp(66781) := x"3082";
    tmp(66782) := x"1841";
    tmp(66783) := x"1041";
    tmp(66784) := x"0821";
    tmp(66785) := x"0820";
    tmp(66786) := x"0820";
    tmp(66787) := x"0820";
    tmp(66788) := x"1020";
    tmp(66789) := x"1020";
    tmp(66790) := x"0820";
    tmp(66791) := x"0820";
    tmp(66792) := x"0820";
    tmp(66793) := x"0020";
    tmp(66794) := x"0020";
    tmp(66795) := x"0820";
    tmp(66796) := x"0840";
    tmp(66797) := x"0840";
    tmp(66798) := x"0840";
    tmp(66799) := x"0840";
    tmp(66800) := x"0820";
    tmp(66801) := x"0820";
    tmp(66802) := x"0820";
    tmp(66803) := x"0841";
    tmp(66804) := x"0841";
    tmp(66805) := x"0860";
    tmp(66806) := x"0860";
    tmp(66807) := x"0040";
    tmp(66808) := x"0020";
    tmp(66809) := x"0040";
    tmp(66810) := x"0840";
    tmp(66811) := x"0820";
    tmp(66812) := x"0820";
    tmp(66813) := x"0820";
    tmp(66814) := x"0820";
    tmp(66815) := x"0820";
    tmp(66816) := x"1820";
    tmp(66817) := x"1820";
    tmp(66818) := x"1820";
    tmp(66819) := x"1820";
    tmp(66820) := x"1820";
    tmp(66821) := x"1000";
    tmp(66822) := x"1820";
    tmp(66823) := x"2020";
    tmp(66824) := x"1820";
    tmp(66825) := x"1000";
    tmp(66826) := x"1000";
    tmp(66827) := x"0800";
    tmp(66828) := x"0800";
    tmp(66829) := x"0800";
    tmp(66830) := x"0800";
    tmp(66831) := x"0800";
    tmp(66832) := x"0800";
    tmp(66833) := x"1000";
    tmp(66834) := x"1800";
    tmp(66835) := x"2000";
    tmp(66836) := x"2800";
    tmp(66837) := x"3000";
    tmp(66838) := x"3800";
    tmp(66839) := x"3800";
    tmp(66840) := x"4000";
    tmp(66841) := x"4000";
    tmp(66842) := x"5000";
    tmp(66843) := x"5800";
    tmp(66844) := x"5800";
    tmp(66845) := x"5800";
    tmp(66846) := x"5800";
    tmp(66847) := x"5820";
    tmp(66848) := x"3000";
    tmp(66849) := x"2800";
    tmp(66850) := x"4000";
    tmp(66851) := x"4800";
    tmp(66852) := x"5000";
    tmp(66853) := x"5800";
    tmp(66854) := x"5800";
    tmp(66855) := x"5800";
    tmp(66856) := x"5800";
    tmp(66857) := x"6000";
    tmp(66858) := x"6800";
    tmp(66859) := x"6020";
    tmp(66860) := x"6020";
    tmp(66861) := x"8020";
    tmp(66862) := x"7020";
    tmp(66863) := x"6820";
    tmp(66864) := x"6820";
    tmp(66865) := x"7020";
    tmp(66866) := x"5820";
    tmp(66867) := x"5000";
    tmp(66868) := x"5800";
    tmp(66869) := x"5800";
    tmp(66870) := x"4800";
    tmp(66871) := x"6000";
    tmp(66872) := x"6800";
    tmp(66873) := x"7000";
    tmp(66874) := x"7000";
    tmp(66875) := x"6800";
    tmp(66876) := x"6000";
    tmp(66877) := x"6000";
    tmp(66878) := x"5800";
    tmp(66879) := x"7000";
    tmp(66880) := x"7820";
    tmp(66881) := x"7820";
    tmp(66882) := x"5000";
    tmp(66883) := x"5820";
    tmp(66884) := x"4861";
    tmp(66885) := x"2861";
    tmp(66886) := x"1861";
    tmp(66887) := x"1061";
    tmp(66888) := x"1061";
    tmp(66889) := x"1061";
    tmp(66890) := x"1061";
    tmp(66891) := x"1061";
    tmp(66892) := x"0841";
    tmp(66893) := x"0841";
    tmp(66894) := x"0840";
    tmp(66895) := x"0840";
    tmp(66896) := x"0840";
    tmp(66897) := x"0840";
    tmp(66898) := x"0840";
    tmp(66899) := x"0841";
    tmp(66900) := x"1061";
    tmp(66901) := x"1081";
    tmp(66902) := x"10a2";
    tmp(66903) := x"18c2";
    tmp(66904) := x"18e3";
    tmp(66905) := x"2104";
    tmp(66906) := x"2125";
    tmp(66907) := x"2946";
    tmp(66908) := x"3187";
    tmp(66909) := x"31a7";
    tmp(66910) := x"39c9";
    tmp(66911) := x"420a";
    tmp(66912) := x"422a";
    tmp(66913) := x"422b";
    tmp(66914) := x"4a4c";
    tmp(66915) := x"524c";
    tmp(66916) := x"526c";
    tmp(66917) := x"528d";
    tmp(66918) := x"5ace";
    tmp(66919) := x"5aaf";
    tmp(66920) := x"5acf";
    tmp(66921) := x"62ef";
    tmp(66922) := x"62f0";
    tmp(66923) := x"6b31";
    tmp(66924) := x"7372";
    tmp(66925) := x"7373";
    tmp(66926) := x"7bb4";
    tmp(66927) := x"8c15";
    tmp(66928) := x"9498";
    tmp(66929) := x"9cb9";
    tmp(66930) := x"a4fb";
    tmp(66931) := x"ad3a";
    tmp(66932) := x"bd7b";
    tmp(66933) := x"c5de";
    tmp(66934) := x"c61f";
    tmp(66935) := x"ce3f";
    tmp(66936) := x"ce5f";
    tmp(66937) := x"ce3f";
    tmp(66938) := x"ce3f";
    tmp(66939) := x"d65f";
    tmp(66940) := x"ce1f";
    tmp(66941) := x"ce1f";
    tmp(66942) := x"c5ff";
    tmp(66943) := x"c5fe";
    tmp(66944) := x"bd9d";
    tmp(66945) := x"bd9d";
    tmp(66946) := x"bdbd";
    tmp(66947) := x"a4f9";
    tmp(66948) := x"ad59";
    tmp(66949) := x"9cd7";
    tmp(66950) := x"9475";
    tmp(66951) := x"8c55";
    tmp(66952) := x"83f3";
    tmp(66953) := x"7bd1";
    tmp(66954) := x"7bb1";
    tmp(66955) := x"7bb1";
    tmp(66956) := x"73b1";
    tmp(66957) := x"6b70";
    tmp(66958) := x"634f";
    tmp(66959) := x"5b0d";
    tmp(66960) := x"0000";
    tmp(66961) := x"0800";
    tmp(66962) := x"0800";
    tmp(66963) := x"0800";
    tmp(66964) := x"0800";
    tmp(66965) := x"0800";
    tmp(66966) := x"0800";
    tmp(66967) := x"0800";
    tmp(66968) := x"0800";
    tmp(66969) := x"0800";
    tmp(66970) := x"0800";
    tmp(66971) := x"0800";
    tmp(66972) := x"0800";
    tmp(66973) := x"0800";
    tmp(66974) := x"1000";
    tmp(66975) := x"1000";
    tmp(66976) := x"0800";
    tmp(66977) := x"0800";
    tmp(66978) := x"0800";
    tmp(66979) := x"0800";
    tmp(66980) := x"0800";
    tmp(66981) := x"0800";
    tmp(66982) := x"1000";
    tmp(66983) := x"1000";
    tmp(66984) := x"0800";
    tmp(66985) := x"1000";
    tmp(66986) := x"0800";
    tmp(66987) := x"0800";
    tmp(66988) := x"0800";
    tmp(66989) := x"0800";
    tmp(66990) := x"0800";
    tmp(66991) := x"1000";
    tmp(66992) := x"1000";
    tmp(66993) := x"1000";
    tmp(66994) := x"1000";
    tmp(66995) := x"1000";
    tmp(66996) := x"0800";
    tmp(66997) := x"0800";
    tmp(66998) := x"0800";
    tmp(66999) := x"1000";
    tmp(67000) := x"1000";
    tmp(67001) := x"1800";
    tmp(67002) := x"2020";
    tmp(67003) := x"2020";
    tmp(67004) := x"2820";
    tmp(67005) := x"2820";
    tmp(67006) := x"2841";
    tmp(67007) := x"3061";
    tmp(67008) := x"3061";
    tmp(67009) := x"2861";
    tmp(67010) := x"3061";
    tmp(67011) := x"2841";
    tmp(67012) := x"2020";
    tmp(67013) := x"1820";
    tmp(67014) := x"1821";
    tmp(67015) := x"1821";
    tmp(67016) := x"1841";
    tmp(67017) := x"1041";
    tmp(67018) := x"0841";
    tmp(67019) := x"0841";
    tmp(67020) := x"1062";
    tmp(67021) := x"1061";
    tmp(67022) := x"0841";
    tmp(67023) := x"0021";
    tmp(67024) := x"0021";
    tmp(67025) := x"0821";
    tmp(67026) := x"0820";
    tmp(67027) := x"0800";
    tmp(67028) := x"0800";
    tmp(67029) := x"0820";
    tmp(67030) := x"0820";
    tmp(67031) := x"0840";
    tmp(67032) := x"0840";
    tmp(67033) := x"0860";
    tmp(67034) := x"0860";
    tmp(67035) := x"0860";
    tmp(67036) := x"0860";
    tmp(67037) := x"0040";
    tmp(67038) := x"0040";
    tmp(67039) := x"0040";
    tmp(67040) := x"0840";
    tmp(67041) := x"0840";
    tmp(67042) := x"0040";
    tmp(67043) := x"0040";
    tmp(67044) := x"0840";
    tmp(67045) := x"0040";
    tmp(67046) := x"0020";
    tmp(67047) := x"0020";
    tmp(67048) := x"0840";
    tmp(67049) := x"0840";
    tmp(67050) := x"0820";
    tmp(67051) := x"0820";
    tmp(67052) := x"0000";
    tmp(67053) := x"0020";
    tmp(67054) := x"0820";
    tmp(67055) := x"0820";
    tmp(67056) := x"0820";
    tmp(67057) := x"1020";
    tmp(67058) := x"1020";
    tmp(67059) := x"1020";
    tmp(67060) := x"1020";
    tmp(67061) := x"1800";
    tmp(67062) := x"2020";
    tmp(67063) := x"2020";
    tmp(67064) := x"1800";
    tmp(67065) := x"1000";
    tmp(67066) := x"1000";
    tmp(67067) := x"0800";
    tmp(67068) := x"0800";
    tmp(67069) := x"0800";
    tmp(67070) := x"0800";
    tmp(67071) := x"0800";
    tmp(67072) := x"1000";
    tmp(67073) := x"1800";
    tmp(67074) := x"1800";
    tmp(67075) := x"2000";
    tmp(67076) := x"2800";
    tmp(67077) := x"3000";
    tmp(67078) := x"3000";
    tmp(67079) := x"3800";
    tmp(67080) := x"4000";
    tmp(67081) := x"4000";
    tmp(67082) := x"4800";
    tmp(67083) := x"5000";
    tmp(67084) := x"5000";
    tmp(67085) := x"5800";
    tmp(67086) := x"5820";
    tmp(67087) := x"4820";
    tmp(67088) := x"2800";
    tmp(67089) := x"3000";
    tmp(67090) := x"4000";
    tmp(67091) := x"4800";
    tmp(67092) := x"5000";
    tmp(67093) := x"5000";
    tmp(67094) := x"5800";
    tmp(67095) := x"5800";
    tmp(67096) := x"5800";
    tmp(67097) := x"6000";
    tmp(67098) := x"5800";
    tmp(67099) := x"5800";
    tmp(67100) := x"7020";
    tmp(67101) := x"7020";
    tmp(67102) := x"6800";
    tmp(67103) := x"6820";
    tmp(67104) := x"7020";
    tmp(67105) := x"6820";
    tmp(67106) := x"5800";
    tmp(67107) := x"5800";
    tmp(67108) := x"6000";
    tmp(67109) := x"5800";
    tmp(67110) := x"5800";
    tmp(67111) := x"5800";
    tmp(67112) := x"6000";
    tmp(67113) := x"6800";
    tmp(67114) := x"6800";
    tmp(67115) := x"6000";
    tmp(67116) := x"6000";
    tmp(67117) := x"5800";
    tmp(67118) := x"6000";
    tmp(67119) := x"7020";
    tmp(67120) := x"8020";
    tmp(67121) := x"5800";
    tmp(67122) := x"3820";
    tmp(67123) := x"3061";
    tmp(67124) := x"2081";
    tmp(67125) := x"1881";
    tmp(67126) := x"1081";
    tmp(67127) := x"1081";
    tmp(67128) := x"1081";
    tmp(67129) := x"1061";
    tmp(67130) := x"1061";
    tmp(67131) := x"1061";
    tmp(67132) := x"1061";
    tmp(67133) := x"0841";
    tmp(67134) := x"0840";
    tmp(67135) := x"0840";
    tmp(67136) := x"0840";
    tmp(67137) := x"0840";
    tmp(67138) := x"0840";
    tmp(67139) := x"0840";
    tmp(67140) := x"0841";
    tmp(67141) := x"1061";
    tmp(67142) := x"1081";
    tmp(67143) := x"10a2";
    tmp(67144) := x"18c3";
    tmp(67145) := x"20e3";
    tmp(67146) := x"2104";
    tmp(67147) := x"2925";
    tmp(67148) := x"2966";
    tmp(67149) := x"3187";
    tmp(67150) := x"39c8";
    tmp(67151) := x"39c9";
    tmp(67152) := x"420a";
    tmp(67153) := x"4a4b";
    tmp(67154) := x"4a2b";
    tmp(67155) := x"4a4c";
    tmp(67156) := x"526d";
    tmp(67157) := x"528d";
    tmp(67158) := x"5ace";
    tmp(67159) := x"5aae";
    tmp(67160) := x"62cf";
    tmp(67161) := x"62ef";
    tmp(67162) := x"62f0";
    tmp(67163) := x"6b31";
    tmp(67164) := x"7372";
    tmp(67165) := x"7b93";
    tmp(67166) := x"8c15";
    tmp(67167) := x"8c36";
    tmp(67168) := x"8c57";
    tmp(67169) := x"9cd9";
    tmp(67170) := x"a4d9";
    tmp(67171) := x"b53c";
    tmp(67172) := x"b53d";
    tmp(67173) := x"bdbf";
    tmp(67174) := x"c63f";
    tmp(67175) := x"ce3f";
    tmp(67176) := x"ce7f";
    tmp(67177) := x"d67f";
    tmp(67178) := x"ce1f";
    tmp(67179) := x"c5ff";
    tmp(67180) := x"ce3f";
    tmp(67181) := x"ce1f";
    tmp(67182) := x"bdde";
    tmp(67183) := x"bdde";
    tmp(67184) := x"b59d";
    tmp(67185) := x"b55b";
    tmp(67186) := x"ad3a";
    tmp(67187) := x"a4f8";
    tmp(67188) := x"9cb7";
    tmp(67189) := x"9497";
    tmp(67190) := x"8c55";
    tmp(67191) := x"8c14";
    tmp(67192) := x"83f3";
    tmp(67193) := x"7bd2";
    tmp(67194) := x"7bd1";
    tmp(67195) := x"6b70";
    tmp(67196) := x"6b50";
    tmp(67197) := x"632f";
    tmp(67198) := x"632e";
    tmp(67199) := x"5acc";
    tmp(67200) := x"0000";
    tmp(67201) := x"0800";
    tmp(67202) := x"0800";
    tmp(67203) := x"0800";
    tmp(67204) := x"0800";
    tmp(67205) := x"0800";
    tmp(67206) := x"0800";
    tmp(67207) := x"0800";
    tmp(67208) := x"0800";
    tmp(67209) := x"0800";
    tmp(67210) := x"0800";
    tmp(67211) := x"0800";
    tmp(67212) := x"0800";
    tmp(67213) := x"0800";
    tmp(67214) := x"0800";
    tmp(67215) := x"0800";
    tmp(67216) := x"0800";
    tmp(67217) := x"0800";
    tmp(67218) := x"0800";
    tmp(67219) := x"0800";
    tmp(67220) := x"0800";
    tmp(67221) := x"0800";
    tmp(67222) := x"0800";
    tmp(67223) := x"0800";
    tmp(67224) := x"0800";
    tmp(67225) := x"0800";
    tmp(67226) := x"0800";
    tmp(67227) := x"0800";
    tmp(67228) := x"0800";
    tmp(67229) := x"0800";
    tmp(67230) := x"0800";
    tmp(67231) := x"0800";
    tmp(67232) := x"0800";
    tmp(67233) := x"0800";
    tmp(67234) := x"0800";
    tmp(67235) := x"0800";
    tmp(67236) := x"1000";
    tmp(67237) := x"1000";
    tmp(67238) := x"1000";
    tmp(67239) := x"1800";
    tmp(67240) := x"1800";
    tmp(67241) := x"1000";
    tmp(67242) := x"1820";
    tmp(67243) := x"2020";
    tmp(67244) := x"2020";
    tmp(67245) := x"2841";
    tmp(67246) := x"2841";
    tmp(67247) := x"2861";
    tmp(67248) := x"2861";
    tmp(67249) := x"2061";
    tmp(67250) := x"1861";
    tmp(67251) := x"1061";
    tmp(67252) := x"0841";
    tmp(67253) := x"0841";
    tmp(67254) := x"0841";
    tmp(67255) := x"0842";
    tmp(67256) := x"0062";
    tmp(67257) := x"0042";
    tmp(67258) := x"0062";
    tmp(67259) := x"0062";
    tmp(67260) := x"0041";
    tmp(67261) := x"0041";
    tmp(67262) := x"0041";
    tmp(67263) := x"0041";
    tmp(67264) := x"0021";
    tmp(67265) := x"0020";
    tmp(67266) := x"0000";
    tmp(67267) := x"0000";
    tmp(67268) := x"0840";
    tmp(67269) := x"0860";
    tmp(67270) := x"0860";
    tmp(67271) := x"0860";
    tmp(67272) := x"0860";
    tmp(67273) := x"0840";
    tmp(67274) := x"0040";
    tmp(67275) := x"0040";
    tmp(67276) := x"0040";
    tmp(67277) := x"0040";
    tmp(67278) := x"0840";
    tmp(67279) := x"0040";
    tmp(67280) := x"0040";
    tmp(67281) := x"0020";
    tmp(67282) := x"0020";
    tmp(67283) := x"0840";
    tmp(67284) := x"0820";
    tmp(67285) := x"0820";
    tmp(67286) := x"0020";
    tmp(67287) := x"0020";
    tmp(67288) := x"0040";
    tmp(67289) := x"0020";
    tmp(67290) := x"0820";
    tmp(67291) := x"0000";
    tmp(67292) := x"0000";
    tmp(67293) := x"0820";
    tmp(67294) := x"0820";
    tmp(67295) := x"0820";
    tmp(67296) := x"0820";
    tmp(67297) := x"0820";
    tmp(67298) := x"0820";
    tmp(67299) := x"0800";
    tmp(67300) := x"1000";
    tmp(67301) := x"2000";
    tmp(67302) := x"2820";
    tmp(67303) := x"2820";
    tmp(67304) := x"2020";
    tmp(67305) := x"1000";
    tmp(67306) := x"1800";
    tmp(67307) := x"1000";
    tmp(67308) := x"0800";
    tmp(67309) := x"0800";
    tmp(67310) := x"1000";
    tmp(67311) := x"1000";
    tmp(67312) := x"1000";
    tmp(67313) := x"1000";
    tmp(67314) := x"1000";
    tmp(67315) := x"1800";
    tmp(67316) := x"2000";
    tmp(67317) := x"2800";
    tmp(67318) := x"3000";
    tmp(67319) := x"3800";
    tmp(67320) := x"4000";
    tmp(67321) := x"4800";
    tmp(67322) := x"4800";
    tmp(67323) := x"5020";
    tmp(67324) := x"5820";
    tmp(67325) := x"5820";
    tmp(67326) := x"5820";
    tmp(67327) := x"3000";
    tmp(67328) := x"2000";
    tmp(67329) := x"3800";
    tmp(67330) := x"4800";
    tmp(67331) := x"5000";
    tmp(67332) := x"5000";
    tmp(67333) := x"5020";
    tmp(67334) := x"6020";
    tmp(67335) := x"5000";
    tmp(67336) := x"5800";
    tmp(67337) := x"5820";
    tmp(67338) := x"5000";
    tmp(67339) := x"6800";
    tmp(67340) := x"6820";
    tmp(67341) := x"6820";
    tmp(67342) := x"6820";
    tmp(67343) := x"6820";
    tmp(67344) := x"6820";
    tmp(67345) := x"6000";
    tmp(67346) := x"6000";
    tmp(67347) := x"6020";
    tmp(67348) := x"6020";
    tmp(67349) := x"5820";
    tmp(67350) := x"5800";
    tmp(67351) := x"5800";
    tmp(67352) := x"6820";
    tmp(67353) := x"6000";
    tmp(67354) := x"6800";
    tmp(67355) := x"6800";
    tmp(67356) := x"6000";
    tmp(67357) := x"6000";
    tmp(67358) := x"6820";
    tmp(67359) := x"7020";
    tmp(67360) := x"6000";
    tmp(67361) := x"3820";
    tmp(67362) := x"2881";
    tmp(67363) := x"1881";
    tmp(67364) := x"1881";
    tmp(67365) := x"1081";
    tmp(67366) := x"1081";
    tmp(67367) := x"1081";
    tmp(67368) := x"1061";
    tmp(67369) := x"1061";
    tmp(67370) := x"1061";
    tmp(67371) := x"1061";
    tmp(67372) := x"1041";
    tmp(67373) := x"0841";
    tmp(67374) := x"0840";
    tmp(67375) := x"0840";
    tmp(67376) := x"0840";
    tmp(67377) := x"0840";
    tmp(67378) := x"0840";
    tmp(67379) := x"0840";
    tmp(67380) := x"0840";
    tmp(67381) := x"0841";
    tmp(67382) := x"1061";
    tmp(67383) := x"1081";
    tmp(67384) := x"18a2";
    tmp(67385) := x"18e3";
    tmp(67386) := x"2104";
    tmp(67387) := x"2925";
    tmp(67388) := x"2945";
    tmp(67389) := x"3166";
    tmp(67390) := x"39a7";
    tmp(67391) := x"39c8";
    tmp(67392) := x"41ea";
    tmp(67393) := x"420a";
    tmp(67394) := x"4a2b";
    tmp(67395) := x"4a4c";
    tmp(67396) := x"526d";
    tmp(67397) := x"528d";
    tmp(67398) := x"528e";
    tmp(67399) := x"5aae";
    tmp(67400) := x"5aae";
    tmp(67401) := x"62cf";
    tmp(67402) := x"6b10";
    tmp(67403) := x"6b52";
    tmp(67404) := x"7352";
    tmp(67405) := x"7373";
    tmp(67406) := x"7bd4";
    tmp(67407) := x"7bf5";
    tmp(67408) := x"9458";
    tmp(67409) := x"a4da";
    tmp(67410) := x"a4fb";
    tmp(67411) := x"b57d";
    tmp(67412) := x"b59e";
    tmp(67413) := x"bdff";
    tmp(67414) := x"c63f";
    tmp(67415) := x"c61f";
    tmp(67416) := x"c5ff";
    tmp(67417) := x"c61f";
    tmp(67418) := x"c61f";
    tmp(67419) := x"c61e";
    tmp(67420) := x"bdde";
    tmp(67421) := x"c5df";
    tmp(67422) := x"c5dd";
    tmp(67423) := x"bd9c";
    tmp(67424) := x"ad3b";
    tmp(67425) := x"a4d9";
    tmp(67426) := x"ad3a";
    tmp(67427) := x"94b7";
    tmp(67428) := x"9497";
    tmp(67429) := x"8c55";
    tmp(67430) := x"83f4";
    tmp(67431) := x"7bd3";
    tmp(67432) := x"7bb1";
    tmp(67433) := x"7391";
    tmp(67434) := x"7390";
    tmp(67435) := x"6b50";
    tmp(67436) := x"6b2f";
    tmp(67437) := x"630e";
    tmp(67438) := x"62ed";
    tmp(67439) := x"5acc";
    tmp(67440) := x"0000";
    tmp(67441) := x"0800";
    tmp(67442) := x"0800";
    tmp(67443) := x"0800";
    tmp(67444) := x"0800";
    tmp(67445) := x"0800";
    tmp(67446) := x"0800";
    tmp(67447) := x"0800";
    tmp(67448) := x"0800";
    tmp(67449) := x"0800";
    tmp(67450) := x"0800";
    tmp(67451) := x"0800";
    tmp(67452) := x"0800";
    tmp(67453) := x"0800";
    tmp(67454) := x"0800";
    tmp(67455) := x"0800";
    tmp(67456) := x"0800";
    tmp(67457) := x"0800";
    tmp(67458) := x"1000";
    tmp(67459) := x"1000";
    tmp(67460) := x"0800";
    tmp(67461) := x"0800";
    tmp(67462) := x"0800";
    tmp(67463) := x"0800";
    tmp(67464) := x"0800";
    tmp(67465) := x"0800";
    tmp(67466) := x"0800";
    tmp(67467) := x"0800";
    tmp(67468) := x"0800";
    tmp(67469) := x"0800";
    tmp(67470) := x"0800";
    tmp(67471) := x"0800";
    tmp(67472) := x"0800";
    tmp(67473) := x"1000";
    tmp(67474) := x"1000";
    tmp(67475) := x"1820";
    tmp(67476) := x"1820";
    tmp(67477) := x"1021";
    tmp(67478) := x"1021";
    tmp(67479) := x"0821";
    tmp(67480) := x"0841";
    tmp(67481) := x"0841";
    tmp(67482) := x"0841";
    tmp(67483) := x"0841";
    tmp(67484) := x"0841";
    tmp(67485) := x"0841";
    tmp(67486) := x"0841";
    tmp(67487) := x"0841";
    tmp(67488) := x"0841";
    tmp(67489) := x"0041";
    tmp(67490) := x"0042";
    tmp(67491) := x"0062";
    tmp(67492) := x"0042";
    tmp(67493) := x"0062";
    tmp(67494) := x"0062";
    tmp(67495) := x"0062";
    tmp(67496) := x"0062";
    tmp(67497) := x"0062";
    tmp(67498) := x"0062";
    tmp(67499) := x"0041";
    tmp(67500) := x"0041";
    tmp(67501) := x"0041";
    tmp(67502) := x"0041";
    tmp(67503) := x"0021";
    tmp(67504) := x"0020";
    tmp(67505) := x"0020";
    tmp(67506) := x"0840";
    tmp(67507) := x"0840";
    tmp(67508) := x"0060";
    tmp(67509) := x"0060";
    tmp(67510) := x"0060";
    tmp(67511) := x"0040";
    tmp(67512) := x"0040";
    tmp(67513) := x"0040";
    tmp(67514) := x"0040";
    tmp(67515) := x"0040";
    tmp(67516) := x"0040";
    tmp(67517) := x"0040";
    tmp(67518) := x"0040";
    tmp(67519) := x"0840";
    tmp(67520) := x"0840";
    tmp(67521) := x"0840";
    tmp(67522) := x"0840";
    tmp(67523) := x"0820";
    tmp(67524) := x"0840";
    tmp(67525) := x"0820";
    tmp(67526) := x"0820";
    tmp(67527) := x"0840";
    tmp(67528) := x"0040";
    tmp(67529) := x"0820";
    tmp(67530) := x"0820";
    tmp(67531) := x"0020";
    tmp(67532) := x"0820";
    tmp(67533) := x"0820";
    tmp(67534) := x"0800";
    tmp(67535) := x"0800";
    tmp(67536) := x"0820";
    tmp(67537) := x"1020";
    tmp(67538) := x"0820";
    tmp(67539) := x"1000";
    tmp(67540) := x"1800";
    tmp(67541) := x"1800";
    tmp(67542) := x"2020";
    tmp(67543) := x"2820";
    tmp(67544) := x"2820";
    tmp(67545) := x"2000";
    tmp(67546) := x"2000";
    tmp(67547) := x"1800";
    tmp(67548) := x"1000";
    tmp(67549) := x"1000";
    tmp(67550) := x"1000";
    tmp(67551) := x"1000";
    tmp(67552) := x"1000";
    tmp(67553) := x"1000";
    tmp(67554) := x"1800";
    tmp(67555) := x"1800";
    tmp(67556) := x"2000";
    tmp(67557) := x"2000";
    tmp(67558) := x"2800";
    tmp(67559) := x"3800";
    tmp(67560) := x"4000";
    tmp(67561) := x"4800";
    tmp(67562) := x"4800";
    tmp(67563) := x"5000";
    tmp(67564) := x"5020";
    tmp(67565) := x"5820";
    tmp(67566) := x"4000";
    tmp(67567) := x"2000";
    tmp(67568) := x"2800";
    tmp(67569) := x"4000";
    tmp(67570) := x"5000";
    tmp(67571) := x"5000";
    tmp(67572) := x"5000";
    tmp(67573) := x"5820";
    tmp(67574) := x"5020";
    tmp(67575) := x"5020";
    tmp(67576) := x"4800";
    tmp(67577) := x"5000";
    tmp(67578) := x"6000";
    tmp(67579) := x"6000";
    tmp(67580) := x"6000";
    tmp(67581) := x"6000";
    tmp(67582) := x"6820";
    tmp(67583) := x"6000";
    tmp(67584) := x"6800";
    tmp(67585) := x"6800";
    tmp(67586) := x"6000";
    tmp(67587) := x"6000";
    tmp(67588) := x"6020";
    tmp(67589) := x"5000";
    tmp(67590) := x"5000";
    tmp(67591) := x"6820";
    tmp(67592) := x"5800";
    tmp(67593) := x"6820";
    tmp(67594) := x"6020";
    tmp(67595) := x"6020";
    tmp(67596) := x"5800";
    tmp(67597) := x"6020";
    tmp(67598) := x"6820";
    tmp(67599) := x"5820";
    tmp(67600) := x"4020";
    tmp(67601) := x"2881";
    tmp(67602) := x"18a1";
    tmp(67603) := x"1881";
    tmp(67604) := x"1881";
    tmp(67605) := x"1881";
    tmp(67606) := x"1081";
    tmp(67607) := x"1081";
    tmp(67608) := x"1061";
    tmp(67609) := x"1061";
    tmp(67610) := x"1061";
    tmp(67611) := x"1061";
    tmp(67612) := x"1041";
    tmp(67613) := x"0841";
    tmp(67614) := x"0840";
    tmp(67615) := x"0840";
    tmp(67616) := x"0840";
    tmp(67617) := x"0840";
    tmp(67618) := x"0840";
    tmp(67619) := x"0840";
    tmp(67620) := x"0840";
    tmp(67621) := x"0841";
    tmp(67622) := x"0841";
    tmp(67623) := x"1061";
    tmp(67624) := x"1081";
    tmp(67625) := x"18a2";
    tmp(67626) := x"18c3";
    tmp(67627) := x"2104";
    tmp(67628) := x"2925";
    tmp(67629) := x"2966";
    tmp(67630) := x"3186";
    tmp(67631) := x"39a8";
    tmp(67632) := x"39c9";
    tmp(67633) := x"420a";
    tmp(67634) := x"422a";
    tmp(67635) := x"4a2b";
    tmp(67636) := x"526c";
    tmp(67637) := x"526d";
    tmp(67638) := x"52ad";
    tmp(67639) := x"5aae";
    tmp(67640) := x"5aae";
    tmp(67641) := x"5acf";
    tmp(67642) := x"62f0";
    tmp(67643) := x"6b51";
    tmp(67644) := x"6b52";
    tmp(67645) := x"7b94";
    tmp(67646) := x"7bb4";
    tmp(67647) := x"8416";
    tmp(67648) := x"8c37";
    tmp(67649) := x"9cdb";
    tmp(67650) := x"ad3b";
    tmp(67651) := x"b59d";
    tmp(67652) := x"bdde";
    tmp(67653) := x"c61f";
    tmp(67654) := x"c5ff";
    tmp(67655) := x"c5fe";
    tmp(67656) := x"c5ff";
    tmp(67657) := x"bdff";
    tmp(67658) := x"bdde";
    tmp(67659) := x"bddd";
    tmp(67660) := x"bdbe";
    tmp(67661) := x"b57c";
    tmp(67662) := x"b55c";
    tmp(67663) := x"ad3b";
    tmp(67664) := x"a4f9";
    tmp(67665) := x"a4d8";
    tmp(67666) := x"a4d7";
    tmp(67667) := x"9475";
    tmp(67668) := x"8c55";
    tmp(67669) := x"8415";
    tmp(67670) := x"83f3";
    tmp(67671) := x"7bb2";
    tmp(67672) := x"7370";
    tmp(67673) := x"6b50";
    tmp(67674) := x"6b50";
    tmp(67675) := x"6b4f";
    tmp(67676) := x"630e";
    tmp(67677) := x"630e";
    tmp(67678) := x"5acd";
    tmp(67679) := x"52cc";
    tmp(67680) := x"0000";
    tmp(67681) := x"0800";
    tmp(67682) := x"0800";
    tmp(67683) := x"0800";
    tmp(67684) := x"0800";
    tmp(67685) := x"0800";
    tmp(67686) := x"0800";
    tmp(67687) := x"0800";
    tmp(67688) := x"0800";
    tmp(67689) := x"0800";
    tmp(67690) := x"0800";
    tmp(67691) := x"0800";
    tmp(67692) := x"0800";
    tmp(67693) := x"0800";
    tmp(67694) := x"0800";
    tmp(67695) := x"0800";
    tmp(67696) := x"1000";
    tmp(67697) := x"1000";
    tmp(67698) := x"1000";
    tmp(67699) := x"0800";
    tmp(67700) := x"0800";
    tmp(67701) := x"0800";
    tmp(67702) := x"0800";
    tmp(67703) := x"0800";
    tmp(67704) := x"0800";
    tmp(67705) := x"0800";
    tmp(67706) := x"0800";
    tmp(67707) := x"0800";
    tmp(67708) := x"0800";
    tmp(67709) := x"1000";
    tmp(67710) := x"1000";
    tmp(67711) := x"1020";
    tmp(67712) := x"1020";
    tmp(67713) := x"0820";
    tmp(67714) := x"0820";
    tmp(67715) := x"0841";
    tmp(67716) := x"0841";
    tmp(67717) := x"0862";
    tmp(67718) := x"0062";
    tmp(67719) := x"0062";
    tmp(67720) := x"0062";
    tmp(67721) := x"0062";
    tmp(67722) := x"0062";
    tmp(67723) := x"0042";
    tmp(67724) := x"0042";
    tmp(67725) := x"0042";
    tmp(67726) := x"0042";
    tmp(67727) := x"0042";
    tmp(67728) := x"0042";
    tmp(67729) := x"0062";
    tmp(67730) := x"0062";
    tmp(67731) := x"0062";
    tmp(67732) := x"0061";
    tmp(67733) := x"0062";
    tmp(67734) := x"0061";
    tmp(67735) := x"0041";
    tmp(67736) := x"0041";
    tmp(67737) := x"0041";
    tmp(67738) := x"0041";
    tmp(67739) := x"0041";
    tmp(67740) := x"0041";
    tmp(67741) := x"0041";
    tmp(67742) := x"0021";
    tmp(67743) := x"0020";
    tmp(67744) := x"0020";
    tmp(67745) := x"0040";
    tmp(67746) := x"0860";
    tmp(67747) := x"0040";
    tmp(67748) := x"0040";
    tmp(67749) := x"0040";
    tmp(67750) := x"0040";
    tmp(67751) := x"0040";
    tmp(67752) := x"0040";
    tmp(67753) := x"0040";
    tmp(67754) := x"0040";
    tmp(67755) := x"0040";
    tmp(67756) := x"0040";
    tmp(67757) := x"0860";
    tmp(67758) := x"0860";
    tmp(67759) := x"0860";
    tmp(67760) := x"0860";
    tmp(67761) := x"0840";
    tmp(67762) := x"0840";
    tmp(67763) := x"0820";
    tmp(67764) := x"0820";
    tmp(67765) := x"0820";
    tmp(67766) := x"0820";
    tmp(67767) := x"0020";
    tmp(67768) := x"0020";
    tmp(67769) := x"0820";
    tmp(67770) := x"0820";
    tmp(67771) := x"0820";
    tmp(67772) := x"0820";
    tmp(67773) := x"0820";
    tmp(67774) := x"1020";
    tmp(67775) := x"1820";
    tmp(67776) := x"1820";
    tmp(67777) := x"1820";
    tmp(67778) := x"1000";
    tmp(67779) := x"1800";
    tmp(67780) := x"2000";
    tmp(67781) := x"2000";
    tmp(67782) := x"1800";
    tmp(67783) := x"2000";
    tmp(67784) := x"2820";
    tmp(67785) := x"2820";
    tmp(67786) := x"2800";
    tmp(67787) := x"1800";
    tmp(67788) := x"1000";
    tmp(67789) := x"1000";
    tmp(67790) := x"1000";
    tmp(67791) := x"1000";
    tmp(67792) := x"0800";
    tmp(67793) := x"1000";
    tmp(67794) := x"1000";
    tmp(67795) := x"1000";
    tmp(67796) := x"1000";
    tmp(67797) := x"1000";
    tmp(67798) := x"2000";
    tmp(67799) := x"3800";
    tmp(67800) := x"4000";
    tmp(67801) := x"4800";
    tmp(67802) := x"4000";
    tmp(67803) := x"4800";
    tmp(67804) := x"4800";
    tmp(67805) := x"4800";
    tmp(67806) := x"2800";
    tmp(67807) := x"1800";
    tmp(67808) := x"3000";
    tmp(67809) := x"4800";
    tmp(67810) := x"5000";
    tmp(67811) := x"5000";
    tmp(67812) := x"5020";
    tmp(67813) := x"5020";
    tmp(67814) := x"4000";
    tmp(67815) := x"4800";
    tmp(67816) := x"4800";
    tmp(67817) := x"5000";
    tmp(67818) := x"6000";
    tmp(67819) := x"6000";
    tmp(67820) := x"6000";
    tmp(67821) := x"6000";
    tmp(67822) := x"5800";
    tmp(67823) := x"5800";
    tmp(67824) := x"6000";
    tmp(67825) := x"6000";
    tmp(67826) := x"5800";
    tmp(67827) := x"5800";
    tmp(67828) := x"5000";
    tmp(67829) := x"5000";
    tmp(67830) := x"6020";
    tmp(67831) := x"6020";
    tmp(67832) := x"6820";
    tmp(67833) := x"6820";
    tmp(67834) := x"6020";
    tmp(67835) := x"5820";
    tmp(67836) := x"5820";
    tmp(67837) := x"6020";
    tmp(67838) := x"5820";
    tmp(67839) := x"4020";
    tmp(67840) := x"2881";
    tmp(67841) := x"20a1";
    tmp(67842) := x"18a1";
    tmp(67843) := x"18a1";
    tmp(67844) := x"1881";
    tmp(67845) := x"1881";
    tmp(67846) := x"1081";
    tmp(67847) := x"1081";
    tmp(67848) := x"1061";
    tmp(67849) := x"1061";
    tmp(67850) := x"1061";
    tmp(67851) := x"1061";
    tmp(67852) := x"0841";
    tmp(67853) := x"0841";
    tmp(67854) := x"0840";
    tmp(67855) := x"0840";
    tmp(67856) := x"0840";
    tmp(67857) := x"0840";
    tmp(67858) := x"0840";
    tmp(67859) := x"0840";
    tmp(67860) := x"0840";
    tmp(67861) := x"0840";
    tmp(67862) := x"0841";
    tmp(67863) := x"0841";
    tmp(67864) := x"1061";
    tmp(67865) := x"1081";
    tmp(67866) := x"18a2";
    tmp(67867) := x"18e3";
    tmp(67868) := x"2104";
    tmp(67869) := x"2945";
    tmp(67870) := x"2966";
    tmp(67871) := x"3187";
    tmp(67872) := x"39c8";
    tmp(67873) := x"41e9";
    tmp(67874) := x"3a09";
    tmp(67875) := x"422b";
    tmp(67876) := x"4a4b";
    tmp(67877) := x"4a6c";
    tmp(67878) := x"528d";
    tmp(67879) := x"52ae";
    tmp(67880) := x"5ace";
    tmp(67881) := x"5ace";
    tmp(67882) := x"5aef";
    tmp(67883) := x"6331";
    tmp(67884) := x"6b52";
    tmp(67885) := x"7372";
    tmp(67886) := x"7bd4";
    tmp(67887) := x"8416";
    tmp(67888) := x"9478";
    tmp(67889) := x"9cd9";
    tmp(67890) := x"acf9";
    tmp(67891) := x"b59c";
    tmp(67892) := x"b59d";
    tmp(67893) := x"bdbd";
    tmp(67894) := x"bdbd";
    tmp(67895) := x"bdde";
    tmp(67896) := x"bdbd";
    tmp(67897) := x"b5bd";
    tmp(67898) := x"b57b";
    tmp(67899) := x"ad3b";
    tmp(67900) := x"bd9c";
    tmp(67901) := x"ad1b";
    tmp(67902) := x"a4d9";
    tmp(67903) := x"a4d8";
    tmp(67904) := x"a4d8";
    tmp(67905) := x"9c96";
    tmp(67906) := x"8c55";
    tmp(67907) := x"8c14";
    tmp(67908) := x"8c14";
    tmp(67909) := x"7bb3";
    tmp(67910) := x"7391";
    tmp(67911) := x"6b51";
    tmp(67912) := x"6b50";
    tmp(67913) := x"6b4f";
    tmp(67914) := x"6b2f";
    tmp(67915) := x"630f";
    tmp(67916) := x"630e";
    tmp(67917) := x"5aee";
    tmp(67918) := x"5acd";
    tmp(67919) := x"528b";
    tmp(67920) := x"0000";
    tmp(67921) := x"0800";
    tmp(67922) := x"0800";
    tmp(67923) := x"0800";
    tmp(67924) := x"0800";
    tmp(67925) := x"0800";
    tmp(67926) := x"0800";
    tmp(67927) := x"0800";
    tmp(67928) := x"0800";
    tmp(67929) := x"0800";
    tmp(67930) := x"0800";
    tmp(67931) := x"0800";
    tmp(67932) := x"0800";
    tmp(67933) := x"0800";
    tmp(67934) := x"0800";
    tmp(67935) := x"0800";
    tmp(67936) := x"0800";
    tmp(67937) := x"0800";
    tmp(67938) := x"0800";
    tmp(67939) := x"0800";
    tmp(67940) := x"0800";
    tmp(67941) := x"0800";
    tmp(67942) := x"0800";
    tmp(67943) := x"0800";
    tmp(67944) := x"0800";
    tmp(67945) := x"0000";
    tmp(67946) := x"0000";
    tmp(67947) := x"0000";
    tmp(67948) := x"0000";
    tmp(67949) := x"0820";
    tmp(67950) := x"0821";
    tmp(67951) := x"0841";
    tmp(67952) := x"0841";
    tmp(67953) := x"0041";
    tmp(67954) := x"0062";
    tmp(67955) := x"0042";
    tmp(67956) := x"0041";
    tmp(67957) := x"0041";
    tmp(67958) := x"0042";
    tmp(67959) := x"0042";
    tmp(67960) := x"0042";
    tmp(67961) := x"0042";
    tmp(67962) := x"0041";
    tmp(67963) := x"0041";
    tmp(67964) := x"0042";
    tmp(67965) := x"0062";
    tmp(67966) := x"0042";
    tmp(67967) := x"0062";
    tmp(67968) := x"0062";
    tmp(67969) := x"0062";
    tmp(67970) := x"0041";
    tmp(67971) := x"0041";
    tmp(67972) := x"0041";
    tmp(67973) := x"0041";
    tmp(67974) := x"0041";
    tmp(67975) := x"0041";
    tmp(67976) := x"0041";
    tmp(67977) := x"0041";
    tmp(67978) := x"0041";
    tmp(67979) := x"0041";
    tmp(67980) := x"0041";
    tmp(67981) := x"0041";
    tmp(67982) := x"0021";
    tmp(67983) := x"0040";
    tmp(67984) := x"0040";
    tmp(67985) := x"0040";
    tmp(67986) := x"0040";
    tmp(67987) := x"0040";
    tmp(67988) := x"0040";
    tmp(67989) := x"0040";
    tmp(67990) := x"0040";
    tmp(67991) := x"0040";
    tmp(67992) := x"0040";
    tmp(67993) := x"0040";
    tmp(67994) := x"0040";
    tmp(67995) := x"0040";
    tmp(67996) := x"0040";
    tmp(67997) := x"0860";
    tmp(67998) := x"0840";
    tmp(67999) := x"0840";
    tmp(68000) := x"0840";
    tmp(68001) := x"0840";
    tmp(68002) := x"0840";
    tmp(68003) := x"0840";
    tmp(68004) := x"0820";
    tmp(68005) := x"0820";
    tmp(68006) := x"0820";
    tmp(68007) := x"0820";
    tmp(68008) := x"0820";
    tmp(68009) := x"0000";
    tmp(68010) := x"0800";
    tmp(68011) := x"0800";
    tmp(68012) := x"0800";
    tmp(68013) := x"0820";
    tmp(68014) := x"1020";
    tmp(68015) := x"1820";
    tmp(68016) := x"2020";
    tmp(68017) := x"1820";
    tmp(68018) := x"1800";
    tmp(68019) := x"1800";
    tmp(68020) := x"2800";
    tmp(68021) := x"2800";
    tmp(68022) := x"2000";
    tmp(68023) := x"2800";
    tmp(68024) := x"2820";
    tmp(68025) := x"2820";
    tmp(68026) := x"2800";
    tmp(68027) := x"2000";
    tmp(68028) := x"1800";
    tmp(68029) := x"1800";
    tmp(68030) := x"1800";
    tmp(68031) := x"1800";
    tmp(68032) := x"1000";
    tmp(68033) := x"1000";
    tmp(68034) := x"1000";
    tmp(68035) := x"0800";
    tmp(68036) := x"0800";
    tmp(68037) := x"1000";
    tmp(68038) := x"2800";
    tmp(68039) := x"3800";
    tmp(68040) := x"4000";
    tmp(68041) := x"4000";
    tmp(68042) := x"4000";
    tmp(68043) := x"4000";
    tmp(68044) := x"4000";
    tmp(68045) := x"3000";
    tmp(68046) := x"2000";
    tmp(68047) := x"2000";
    tmp(68048) := x"3800";
    tmp(68049) := x"4000";
    tmp(68050) := x"4800";
    tmp(68051) := x"4800";
    tmp(68052) := x"4820";
    tmp(68053) := x"4000";
    tmp(68054) := x"4000";
    tmp(68055) := x"4800";
    tmp(68056) := x"4800";
    tmp(68057) := x"5800";
    tmp(68058) := x"6000";
    tmp(68059) := x"6000";
    tmp(68060) := x"6800";
    tmp(68061) := x"6000";
    tmp(68062) := x"5800";
    tmp(68063) := x"5800";
    tmp(68064) := x"6000";
    tmp(68065) := x"5800";
    tmp(68066) := x"5000";
    tmp(68067) := x"5800";
    tmp(68068) := x"5000";
    tmp(68069) := x"5800";
    tmp(68070) := x"6820";
    tmp(68071) := x"6020";
    tmp(68072) := x"7020";
    tmp(68073) := x"5820";
    tmp(68074) := x"4820";
    tmp(68075) := x"5020";
    tmp(68076) := x"4820";
    tmp(68077) := x"5041";
    tmp(68078) := x"3861";
    tmp(68079) := x"28a1";
    tmp(68080) := x"20c2";
    tmp(68081) := x"18a2";
    tmp(68082) := x"18a2";
    tmp(68083) := x"18a1";
    tmp(68084) := x"1881";
    tmp(68085) := x"1881";
    tmp(68086) := x"1081";
    tmp(68087) := x"1081";
    tmp(68088) := x"1061";
    tmp(68089) := x"1061";
    tmp(68090) := x"1061";
    tmp(68091) := x"1061";
    tmp(68092) := x"0841";
    tmp(68093) := x"0841";
    tmp(68094) := x"0840";
    tmp(68095) := x"0840";
    tmp(68096) := x"0840";
    tmp(68097) := x"0840";
    tmp(68098) := x"0840";
    tmp(68099) := x"0840";
    tmp(68100) := x"0820";
    tmp(68101) := x"0820";
    tmp(68102) := x"0840";
    tmp(68103) := x"0841";
    tmp(68104) := x"0861";
    tmp(68105) := x"1061";
    tmp(68106) := x"1081";
    tmp(68107) := x"18a2";
    tmp(68108) := x"18e3";
    tmp(68109) := x"2104";
    tmp(68110) := x"2945";
    tmp(68111) := x"2966";
    tmp(68112) := x"3187";
    tmp(68113) := x"39a8";
    tmp(68114) := x"39e9";
    tmp(68115) := x"420a";
    tmp(68116) := x"420a";
    tmp(68117) := x"422b";
    tmp(68118) := x"4a4b";
    tmp(68119) := x"4a4c";
    tmp(68120) := x"526c";
    tmp(68121) := x"5aad";
    tmp(68122) := x"5ace";
    tmp(68123) := x"62ef";
    tmp(68124) := x"6b30";
    tmp(68125) := x"6b51";
    tmp(68126) := x"7b92";
    tmp(68127) := x"7bf4";
    tmp(68128) := x"8c35";
    tmp(68129) := x"9497";
    tmp(68130) := x"9cd8";
    tmp(68131) := x"a4f9";
    tmp(68132) := x"ad3b";
    tmp(68133) := x"b57c";
    tmp(68134) := x"b57d";
    tmp(68135) := x"ad5c";
    tmp(68136) := x"b55b";
    tmp(68137) := x"ad5b";
    tmp(68138) := x"a53a";
    tmp(68139) := x"a519";
    tmp(68140) := x"a4f9";
    tmp(68141) := x"a4d8";
    tmp(68142) := x"9c76";
    tmp(68143) := x"9c97";
    tmp(68144) := x"9475";
    tmp(68145) := x"8c35";
    tmp(68146) := x"83f4";
    tmp(68147) := x"83d2";
    tmp(68148) := x"7b92";
    tmp(68149) := x"7b92";
    tmp(68150) := x"7371";
    tmp(68151) := x"6b50";
    tmp(68152) := x"6b2f";
    tmp(68153) := x"6b2f";
    tmp(68154) := x"630e";
    tmp(68155) := x"62ee";
    tmp(68156) := x"62ee";
    tmp(68157) := x"5acd";
    tmp(68158) := x"52ac";
    tmp(68159) := x"4a6b";
    tmp(68160) := x"0000";
    tmp(68161) := x"0800";
    tmp(68162) := x"0800";
    tmp(68163) := x"0800";
    tmp(68164) := x"0800";
    tmp(68165) := x"0800";
    tmp(68166) := x"0800";
    tmp(68167) := x"0800";
    tmp(68168) := x"0800";
    tmp(68169) := x"0800";
    tmp(68170) := x"0800";
    tmp(68171) := x"0800";
    tmp(68172) := x"0800";
    tmp(68173) := x"0800";
    tmp(68174) := x"0800";
    tmp(68175) := x"0800";
    tmp(68176) := x"0800";
    tmp(68177) := x"0800";
    tmp(68178) := x"0800";
    tmp(68179) := x"0800";
    tmp(68180) := x"0800";
    tmp(68181) := x"0800";
    tmp(68182) := x"0800";
    tmp(68183) := x"0800";
    tmp(68184) := x"0800";
    tmp(68185) := x"0000";
    tmp(68186) := x"0020";
    tmp(68187) := x"0021";
    tmp(68188) := x"0041";
    tmp(68189) := x"0041";
    tmp(68190) := x"0041";
    tmp(68191) := x"0021";
    tmp(68192) := x"0041";
    tmp(68193) := x"0041";
    tmp(68194) := x"0041";
    tmp(68195) := x"0041";
    tmp(68196) := x"0041";
    tmp(68197) := x"0041";
    tmp(68198) := x"0041";
    tmp(68199) := x"0041";
    tmp(68200) := x"0042";
    tmp(68201) := x"0041";
    tmp(68202) := x"0041";
    tmp(68203) := x"0041";
    tmp(68204) := x"0041";
    tmp(68205) := x"0041";
    tmp(68206) := x"0041";
    tmp(68207) := x"0041";
    tmp(68208) := x"0041";
    tmp(68209) := x"0041";
    tmp(68210) := x"0041";
    tmp(68211) := x"0041";
    tmp(68212) := x"0041";
    tmp(68213) := x"0041";
    tmp(68214) := x"0041";
    tmp(68215) := x"0041";
    tmp(68216) := x"0041";
    tmp(68217) := x"0041";
    tmp(68218) := x"0041";
    tmp(68219) := x"0041";
    tmp(68220) := x"0041";
    tmp(68221) := x"0041";
    tmp(68222) := x"0041";
    tmp(68223) := x"0020";
    tmp(68224) := x"0020";
    tmp(68225) := x"0020";
    tmp(68226) := x"0040";
    tmp(68227) := x"0040";
    tmp(68228) := x"0040";
    tmp(68229) := x"0040";
    tmp(68230) := x"0040";
    tmp(68231) := x"0040";
    tmp(68232) := x"0040";
    tmp(68233) := x"0840";
    tmp(68234) := x"0040";
    tmp(68235) := x"0040";
    tmp(68236) := x"0040";
    tmp(68237) := x"0840";
    tmp(68238) := x"0840";
    tmp(68239) := x"0840";
    tmp(68240) := x"0840";
    tmp(68241) := x"0840";
    tmp(68242) := x"0840";
    tmp(68243) := x"0840";
    tmp(68244) := x"0840";
    tmp(68245) := x"0820";
    tmp(68246) := x"0820";
    tmp(68247) := x"0820";
    tmp(68248) := x"0820";
    tmp(68249) := x"0800";
    tmp(68250) := x"0800";
    tmp(68251) := x"0820";
    tmp(68252) := x"1020";
    tmp(68253) := x"1020";
    tmp(68254) := x"1020";
    tmp(68255) := x"1820";
    tmp(68256) := x"1820";
    tmp(68257) := x"1020";
    tmp(68258) := x"1000";
    tmp(68259) := x"2000";
    tmp(68260) := x"2800";
    tmp(68261) := x"2800";
    tmp(68262) := x"2800";
    tmp(68263) := x"3000";
    tmp(68264) := x"2800";
    tmp(68265) := x"2800";
    tmp(68266) := x"2800";
    tmp(68267) := x"2000";
    tmp(68268) := x"2000";
    tmp(68269) := x"2000";
    tmp(68270) := x"2800";
    tmp(68271) := x"2000";
    tmp(68272) := x"2000";
    tmp(68273) := x"1000";
    tmp(68274) := x"1000";
    tmp(68275) := x"0800";
    tmp(68276) := x"0800";
    tmp(68277) := x"2000";
    tmp(68278) := x"2800";
    tmp(68279) := x"3000";
    tmp(68280) := x"3000";
    tmp(68281) := x"3800";
    tmp(68282) := x"4000";
    tmp(68283) := x"4000";
    tmp(68284) := x"3800";
    tmp(68285) := x"2800";
    tmp(68286) := x"2000";
    tmp(68287) := x"2800";
    tmp(68288) := x"3800";
    tmp(68289) := x"3800";
    tmp(68290) := x"3800";
    tmp(68291) := x"3800";
    tmp(68292) := x"3800";
    tmp(68293) := x"3000";
    tmp(68294) := x"4800";
    tmp(68295) := x"4800";
    tmp(68296) := x"5020";
    tmp(68297) := x"6020";
    tmp(68298) := x"5800";
    tmp(68299) := x"5800";
    tmp(68300) := x"6000";
    tmp(68301) := x"5000";
    tmp(68302) := x"5000";
    tmp(68303) := x"5800";
    tmp(68304) := x"5800";
    tmp(68305) := x"5800";
    tmp(68306) := x"3800";
    tmp(68307) := x"5000";
    tmp(68308) := x"5800";
    tmp(68309) := x"6020";
    tmp(68310) := x"5800";
    tmp(68311) := x"7820";
    tmp(68312) := x"6020";
    tmp(68313) := x"4840";
    tmp(68314) := x"4820";
    tmp(68315) := x"3820";
    tmp(68316) := x"4061";
    tmp(68317) := x"3881";
    tmp(68318) := x"28c2";
    tmp(68319) := x"20c2";
    tmp(68320) := x"18a2";
    tmp(68321) := x"18a2";
    tmp(68322) := x"18a1";
    tmp(68323) := x"18a1";
    tmp(68324) := x"1881";
    tmp(68325) := x"1081";
    tmp(68326) := x"1081";
    tmp(68327) := x"1081";
    tmp(68328) := x"1061";
    tmp(68329) := x"1061";
    tmp(68330) := x"1061";
    tmp(68331) := x"1061";
    tmp(68332) := x"0840";
    tmp(68333) := x"0840";
    tmp(68334) := x"0840";
    tmp(68335) := x"0840";
    tmp(68336) := x"0840";
    tmp(68337) := x"0840";
    tmp(68338) := x"0840";
    tmp(68339) := x"0840";
    tmp(68340) := x"0820";
    tmp(68341) := x"0820";
    tmp(68342) := x"0840";
    tmp(68343) := x"0840";
    tmp(68344) := x"0841";
    tmp(68345) := x"0861";
    tmp(68346) := x"1061";
    tmp(68347) := x"1081";
    tmp(68348) := x"18a2";
    tmp(68349) := x"18e3";
    tmp(68350) := x"2104";
    tmp(68351) := x"2125";
    tmp(68352) := x"2966";
    tmp(68353) := x"31a7";
    tmp(68354) := x"39a7";
    tmp(68355) := x"39c8";
    tmp(68356) := x"39c9";
    tmp(68357) := x"39e9";
    tmp(68358) := x"420a";
    tmp(68359) := x"420a";
    tmp(68360) := x"422a";
    tmp(68361) := x"4a4b";
    tmp(68362) := x"528c";
    tmp(68363) := x"5aad";
    tmp(68364) := x"5ace";
    tmp(68365) := x"630f";
    tmp(68366) := x"6b50";
    tmp(68367) := x"7371";
    tmp(68368) := x"7bd3";
    tmp(68369) := x"8414";
    tmp(68370) := x"8c75";
    tmp(68371) := x"9497";
    tmp(68372) := x"9cd9";
    tmp(68373) := x"a4fb";
    tmp(68374) := x"a4fb";
    tmp(68375) := x"ad1a";
    tmp(68376) := x"acfa";
    tmp(68377) := x"a4f9";
    tmp(68378) := x"9cf8";
    tmp(68379) := x"9cd7";
    tmp(68380) := x"9496";
    tmp(68381) := x"9476";
    tmp(68382) := x"9455";
    tmp(68383) := x"8c14";
    tmp(68384) := x"8bf3";
    tmp(68385) := x"83d3";
    tmp(68386) := x"7392";
    tmp(68387) := x"7391";
    tmp(68388) := x"7391";
    tmp(68389) := x"7371";
    tmp(68390) := x"6b50";
    tmp(68391) := x"6b2f";
    tmp(68392) := x"632f";
    tmp(68393) := x"632f";
    tmp(68394) := x"62ee";
    tmp(68395) := x"5ace";
    tmp(68396) := x"5aad";
    tmp(68397) := x"528c";
    tmp(68398) := x"526b";
    tmp(68399) := x"4a6b";
    tmp(68400) := x"0000";
    tmp(68401) := x"0800";
    tmp(68402) := x"0800";
    tmp(68403) := x"0020";
    tmp(68404) := x"0020";
    tmp(68405) := x"0020";
    tmp(68406) := x"0021";
    tmp(68407) := x"0021";
    tmp(68408) := x"0021";
    tmp(68409) := x"0021";
    tmp(68410) := x"0021";
    tmp(68411) := x"0041";
    tmp(68412) := x"0021";
    tmp(68413) := x"0021";
    tmp(68414) := x"0021";
    tmp(68415) := x"0020";
    tmp(68416) := x"0020";
    tmp(68417) := x"0020";
    tmp(68418) := x"0020";
    tmp(68419) := x"0000";
    tmp(68420) := x"0020";
    tmp(68421) := x"0020";
    tmp(68422) := x"0020";
    tmp(68423) := x"0021";
    tmp(68424) := x"0041";
    tmp(68425) := x"0041";
    tmp(68426) := x"0041";
    tmp(68427) := x"0021";
    tmp(68428) := x"0021";
    tmp(68429) := x"0021";
    tmp(68430) := x"0021";
    tmp(68431) := x"0021";
    tmp(68432) := x"0021";
    tmp(68433) := x"0021";
    tmp(68434) := x"0021";
    tmp(68435) := x"0041";
    tmp(68436) := x"0041";
    tmp(68437) := x"0041";
    tmp(68438) := x"0041";
    tmp(68439) := x"0041";
    tmp(68440) := x"0041";
    tmp(68441) := x"0041";
    tmp(68442) := x"0041";
    tmp(68443) := x"0041";
    tmp(68444) := x"0041";
    tmp(68445) := x"0041";
    tmp(68446) := x"0041";
    tmp(68447) := x"0041";
    tmp(68448) := x"0041";
    tmp(68449) := x"0041";
    tmp(68450) := x"0041";
    tmp(68451) := x"0041";
    tmp(68452) := x"0041";
    tmp(68453) := x"0041";
    tmp(68454) := x"0041";
    tmp(68455) := x"0041";
    tmp(68456) := x"0041";
    tmp(68457) := x"0061";
    tmp(68458) := x"0041";
    tmp(68459) := x"0041";
    tmp(68460) := x"0041";
    tmp(68461) := x"0041";
    tmp(68462) := x"0021";
    tmp(68463) := x"0020";
    tmp(68464) := x"0020";
    tmp(68465) := x"0020";
    tmp(68466) := x"0020";
    tmp(68467) := x"0040";
    tmp(68468) := x"0040";
    tmp(68469) := x"0040";
    tmp(68470) := x"0040";
    tmp(68471) := x"0060";
    tmp(68472) := x"0040";
    tmp(68473) := x"0040";
    tmp(68474) := x"0040";
    tmp(68475) := x"0020";
    tmp(68476) := x"0040";
    tmp(68477) := x"0040";
    tmp(68478) := x"0840";
    tmp(68479) := x"0840";
    tmp(68480) := x"0840";
    tmp(68481) := x"0840";
    tmp(68482) := x"0840";
    tmp(68483) := x"0840";
    tmp(68484) := x"0840";
    tmp(68485) := x"0820";
    tmp(68486) := x"0820";
    tmp(68487) := x"0800";
    tmp(68488) := x"0800";
    tmp(68489) := x"0820";
    tmp(68490) := x"0820";
    tmp(68491) := x"0820";
    tmp(68492) := x"1020";
    tmp(68493) := x"1020";
    tmp(68494) := x"1820";
    tmp(68495) := x"1020";
    tmp(68496) := x"1020";
    tmp(68497) := x"0800";
    tmp(68498) := x"1000";
    tmp(68499) := x"2000";
    tmp(68500) := x"2800";
    tmp(68501) := x"2800";
    tmp(68502) := x"2800";
    tmp(68503) := x"3000";
    tmp(68504) := x"3020";
    tmp(68505) := x"2800";
    tmp(68506) := x"2800";
    tmp(68507) := x"2800";
    tmp(68508) := x"2800";
    tmp(68509) := x"2800";
    tmp(68510) := x"3000";
    tmp(68511) := x"3000";
    tmp(68512) := x"2820";
    tmp(68513) := x"1820";
    tmp(68514) := x"1000";
    tmp(68515) := x"1000";
    tmp(68516) := x"1000";
    tmp(68517) := x"1800";
    tmp(68518) := x"2000";
    tmp(68519) := x"2000";
    tmp(68520) := x"2800";
    tmp(68521) := x"3800";
    tmp(68522) := x"3800";
    tmp(68523) := x"3800";
    tmp(68524) := x"2800";
    tmp(68525) := x"2000";
    tmp(68526) := x"2000";
    tmp(68527) := x"2800";
    tmp(68528) := x"3000";
    tmp(68529) := x"3000";
    tmp(68530) := x"3000";
    tmp(68531) := x"3000";
    tmp(68532) := x"3000";
    tmp(68533) := x"3800";
    tmp(68534) := x"3800";
    tmp(68535) := x"4800";
    tmp(68536) := x"5820";
    tmp(68537) := x"5820";
    tmp(68538) := x"5800";
    tmp(68539) := x"5000";
    tmp(68540) := x"5000";
    tmp(68541) := x"5000";
    tmp(68542) := x"5000";
    tmp(68543) := x"5000";
    tmp(68544) := x"5000";
    tmp(68545) := x"4000";
    tmp(68546) := x"3800";
    tmp(68547) := x"4800";
    tmp(68548) := x"5820";
    tmp(68549) := x"5800";
    tmp(68550) := x"6820";
    tmp(68551) := x"7020";
    tmp(68552) := x"4040";
    tmp(68553) := x"4061";
    tmp(68554) := x"3840";
    tmp(68555) := x"2861";
    tmp(68556) := x"30a2";
    tmp(68557) := x"28a2";
    tmp(68558) := x"20c2";
    tmp(68559) := x"18a2";
    tmp(68560) := x"18a2";
    tmp(68561) := x"18a2";
    tmp(68562) := x"18a1";
    tmp(68563) := x"18a1";
    tmp(68564) := x"1881";
    tmp(68565) := x"1081";
    tmp(68566) := x"1081";
    tmp(68567) := x"1081";
    tmp(68568) := x"1061";
    tmp(68569) := x"1061";
    tmp(68570) := x"1061";
    tmp(68571) := x"1061";
    tmp(68572) := x"0840";
    tmp(68573) := x"0840";
    tmp(68574) := x"0840";
    tmp(68575) := x"0840";
    tmp(68576) := x"0840";
    tmp(68577) := x"0840";
    tmp(68578) := x"0840";
    tmp(68579) := x"0840";
    tmp(68580) := x"0820";
    tmp(68581) := x"0820";
    tmp(68582) := x"0820";
    tmp(68583) := x"0840";
    tmp(68584) := x"0840";
    tmp(68585) := x"0841";
    tmp(68586) := x"0861";
    tmp(68587) := x"1061";
    tmp(68588) := x"1081";
    tmp(68589) := x"18a2";
    tmp(68590) := x"18c3";
    tmp(68591) := x"2104";
    tmp(68592) := x"2124";
    tmp(68593) := x"2965";
    tmp(68594) := x"3186";
    tmp(68595) := x"3187";
    tmp(68596) := x"3187";
    tmp(68597) := x"31a8";
    tmp(68598) := x"39c8";
    tmp(68599) := x"39c8";
    tmp(68600) := x"39e8";
    tmp(68601) := x"420a";
    tmp(68602) := x"4a2a";
    tmp(68603) := x"4a4b";
    tmp(68604) := x"526c";
    tmp(68605) := x"52cd";
    tmp(68606) := x"5aee";
    tmp(68607) := x"632f";
    tmp(68608) := x"6b50";
    tmp(68609) := x"7bb2";
    tmp(68610) := x"7c13";
    tmp(68611) := x"8c55";
    tmp(68612) := x"9497";
    tmp(68613) := x"9498";
    tmp(68614) := x"9498";
    tmp(68615) := x"9c98";
    tmp(68616) := x"9497";
    tmp(68617) := x"9cb7";
    tmp(68618) := x"9475";
    tmp(68619) := x"9455";
    tmp(68620) := x"8c35";
    tmp(68621) := x"8bf4";
    tmp(68622) := x"83f3";
    tmp(68623) := x"83b3";
    tmp(68624) := x"7bb2";
    tmp(68625) := x"7391";
    tmp(68626) := x"7370";
    tmp(68627) := x"6b50";
    tmp(68628) := x"6b50";
    tmp(68629) := x"6b4f";
    tmp(68630) := x"6b2f";
    tmp(68631) := x"630f";
    tmp(68632) := x"62ee";
    tmp(68633) := x"5aee";
    tmp(68634) := x"5ace";
    tmp(68635) := x"5acd";
    tmp(68636) := x"528d";
    tmp(68637) := x"5aad";
    tmp(68638) := x"4a6a";
    tmp(68639) := x"4a4a";
    tmp(68640) := x"0000";
    tmp(68641) := x"0021";
    tmp(68642) := x"0021";
    tmp(68643) := x"0041";
    tmp(68644) := x"0041";
    tmp(68645) := x"0041";
    tmp(68646) := x"0041";
    tmp(68647) := x"0041";
    tmp(68648) := x"0041";
    tmp(68649) := x"0041";
    tmp(68650) := x"0041";
    tmp(68651) := x"0041";
    tmp(68652) := x"0041";
    tmp(68653) := x"0041";
    tmp(68654) := x"0041";
    tmp(68655) := x"0041";
    tmp(68656) := x"0041";
    tmp(68657) := x"0041";
    tmp(68658) := x"0041";
    tmp(68659) := x"0041";
    tmp(68660) := x"0041";
    tmp(68661) := x"0041";
    tmp(68662) := x"0041";
    tmp(68663) := x"0041";
    tmp(68664) := x"0061";
    tmp(68665) := x"0041";
    tmp(68666) := x"0041";
    tmp(68667) := x"0041";
    tmp(68668) := x"0041";
    tmp(68669) := x"0061";
    tmp(68670) := x"0062";
    tmp(68671) := x"0062";
    tmp(68672) := x"0062";
    tmp(68673) := x"0062";
    tmp(68674) := x"0062";
    tmp(68675) := x"0062";
    tmp(68676) := x"0061";
    tmp(68677) := x"0041";
    tmp(68678) := x"0041";
    tmp(68679) := x"0041";
    tmp(68680) := x"0021";
    tmp(68681) := x"0041";
    tmp(68682) := x"0041";
    tmp(68683) := x"0041";
    tmp(68684) := x"0041";
    tmp(68685) := x"0041";
    tmp(68686) := x"0041";
    tmp(68687) := x"0041";
    tmp(68688) := x"0041";
    tmp(68689) := x"0041";
    tmp(68690) := x"0041";
    tmp(68691) := x"0061";
    tmp(68692) := x"0062";
    tmp(68693) := x"0062";
    tmp(68694) := x"0062";
    tmp(68695) := x"0061";
    tmp(68696) := x"0041";
    tmp(68697) := x"0041";
    tmp(68698) := x"0061";
    tmp(68699) := x"0041";
    tmp(68700) := x"0061";
    tmp(68701) := x"0061";
    tmp(68702) := x"0041";
    tmp(68703) := x"0040";
    tmp(68704) := x"0040";
    tmp(68705) := x"0040";
    tmp(68706) := x"0040";
    tmp(68707) := x"0040";
    tmp(68708) := x"0040";
    tmp(68709) := x"0040";
    tmp(68710) := x"0840";
    tmp(68711) := x"0860";
    tmp(68712) := x"0840";
    tmp(68713) := x"0040";
    tmp(68714) := x"0020";
    tmp(68715) := x"0040";
    tmp(68716) := x"0040";
    tmp(68717) := x"0040";
    tmp(68718) := x"0020";
    tmp(68719) := x"0840";
    tmp(68720) := x"0840";
    tmp(68721) := x"0840";
    tmp(68722) := x"0840";
    tmp(68723) := x"0840";
    tmp(68724) := x"0840";
    tmp(68725) := x"0840";
    tmp(68726) := x"0820";
    tmp(68727) := x"0800";
    tmp(68728) := x"0820";
    tmp(68729) := x"0820";
    tmp(68730) := x"0820";
    tmp(68731) := x"0820";
    tmp(68732) := x"0820";
    tmp(68733) := x"1020";
    tmp(68734) := x"1820";
    tmp(68735) := x"1020";
    tmp(68736) := x"0800";
    tmp(68737) := x"1000";
    tmp(68738) := x"1000";
    tmp(68739) := x"2000";
    tmp(68740) := x"2800";
    tmp(68741) := x"2800";
    tmp(68742) := x"2800";
    tmp(68743) := x"3800";
    tmp(68744) := x"3820";
    tmp(68745) := x"3000";
    tmp(68746) := x"2800";
    tmp(68747) := x"3000";
    tmp(68748) := x"2800";
    tmp(68749) := x"3000";
    tmp(68750) := x"3020";
    tmp(68751) := x"3000";
    tmp(68752) := x"2820";
    tmp(68753) := x"1820";
    tmp(68754) := x"1000";
    tmp(68755) := x"1000";
    tmp(68756) := x"1800";
    tmp(68757) := x"1800";
    tmp(68758) := x"1800";
    tmp(68759) := x"2800";
    tmp(68760) := x"3000";
    tmp(68761) := x"3000";
    tmp(68762) := x"3800";
    tmp(68763) := x"3000";
    tmp(68764) := x"2000";
    tmp(68765) := x"1800";
    tmp(68766) := x"2000";
    tmp(68767) := x"2800";
    tmp(68768) := x"2800";
    tmp(68769) := x"2800";
    tmp(68770) := x"2800";
    tmp(68771) := x"3000";
    tmp(68772) := x"3000";
    tmp(68773) := x"3800";
    tmp(68774) := x"3800";
    tmp(68775) := x"4800";
    tmp(68776) := x"5000";
    tmp(68777) := x"4800";
    tmp(68778) := x"4800";
    tmp(68779) := x"4800";
    tmp(68780) := x"4800";
    tmp(68781) := x"4800";
    tmp(68782) := x"4800";
    tmp(68783) := x"4800";
    tmp(68784) := x"4800";
    tmp(68785) := x"3800";
    tmp(68786) := x"4000";
    tmp(68787) := x"5820";
    tmp(68788) := x"5800";
    tmp(68789) := x"6820";
    tmp(68790) := x"6820";
    tmp(68791) := x"4840";
    tmp(68792) := x"3861";
    tmp(68793) := x"3040";
    tmp(68794) := x"2061";
    tmp(68795) := x"20c2";
    tmp(68796) := x"20a2";
    tmp(68797) := x"20c2";
    tmp(68798) := x"18a2";
    tmp(68799) := x"18a2";
    tmp(68800) := x"18a2";
    tmp(68801) := x"18a2";
    tmp(68802) := x"18a1";
    tmp(68803) := x"18a1";
    tmp(68804) := x"1081";
    tmp(68805) := x"1081";
    tmp(68806) := x"1081";
    tmp(68807) := x"1061";
    tmp(68808) := x"1061";
    tmp(68809) := x"1061";
    tmp(68810) := x"1061";
    tmp(68811) := x"1041";
    tmp(68812) := x"0840";
    tmp(68813) := x"0840";
    tmp(68814) := x"0840";
    tmp(68815) := x"0840";
    tmp(68816) := x"0840";
    tmp(68817) := x"0840";
    tmp(68818) := x"0840";
    tmp(68819) := x"0840";
    tmp(68820) := x"0820";
    tmp(68821) := x"0820";
    tmp(68822) := x"0820";
    tmp(68823) := x"0820";
    tmp(68824) := x"0840";
    tmp(68825) := x"0840";
    tmp(68826) := x"0841";
    tmp(68827) := x"0861";
    tmp(68828) := x"1081";
    tmp(68829) := x"1081";
    tmp(68830) := x"18a2";
    tmp(68831) := x"18e3";
    tmp(68832) := x"2103";
    tmp(68833) := x"2124";
    tmp(68834) := x"2125";
    tmp(68835) := x"2945";
    tmp(68836) := x"2966";
    tmp(68837) := x"2986";
    tmp(68838) := x"3186";
    tmp(68839) := x"3186";
    tmp(68840) := x"31a7";
    tmp(68841) := x"39c8";
    tmp(68842) := x"39e8";
    tmp(68843) := x"4209";
    tmp(68844) := x"4a2a";
    tmp(68845) := x"4a6a";
    tmp(68846) := x"528c";
    tmp(68847) := x"5acd";
    tmp(68848) := x"62ee";
    tmp(68849) := x"6b2f";
    tmp(68850) := x"7391";
    tmp(68851) := x"83f3";
    tmp(68852) := x"8c34";
    tmp(68853) := x"8c54";
    tmp(68854) := x"8c35";
    tmp(68855) := x"8c56";
    tmp(68856) := x"8c55";
    tmp(68857) := x"8c34";
    tmp(68858) := x"8c14";
    tmp(68859) := x"8bf3";
    tmp(68860) := x"83d3";
    tmp(68861) := x"7bb3";
    tmp(68862) := x"7392";
    tmp(68863) := x"7371";
    tmp(68864) := x"7350";
    tmp(68865) := x"7370";
    tmp(68866) := x"6b50";
    tmp(68867) := x"6b4f";
    tmp(68868) := x"6b0f";
    tmp(68869) := x"630f";
    tmp(68870) := x"630f";
    tmp(68871) := x"62ee";
    tmp(68872) := x"62ee";
    tmp(68873) := x"5acd";
    tmp(68874) := x"5acd";
    tmp(68875) := x"5aad";
    tmp(68876) := x"528c";
    tmp(68877) := x"528b";
    tmp(68878) := x"4a4a";
    tmp(68879) := x"422a";
    tmp(68880) := x"0000";
    tmp(68881) := x"0041";
    tmp(68882) := x"0041";
    tmp(68883) := x"0041";
    tmp(68884) := x"0041";
    tmp(68885) := x"0041";
    tmp(68886) := x"0041";
    tmp(68887) := x"0041";
    tmp(68888) := x"0041";
    tmp(68889) := x"0041";
    tmp(68890) := x"0041";
    tmp(68891) := x"0041";
    tmp(68892) := x"0041";
    tmp(68893) := x"0041";
    tmp(68894) := x"0041";
    tmp(68895) := x"0041";
    tmp(68896) := x"0041";
    tmp(68897) := x"0041";
    tmp(68898) := x"0041";
    tmp(68899) := x"0041";
    tmp(68900) := x"0041";
    tmp(68901) := x"0041";
    tmp(68902) := x"0041";
    tmp(68903) := x"0041";
    tmp(68904) := x"0041";
    tmp(68905) := x"0041";
    tmp(68906) := x"0041";
    tmp(68907) := x"0061";
    tmp(68908) := x"0061";
    tmp(68909) := x"0061";
    tmp(68910) := x"0062";
    tmp(68911) := x"0062";
    tmp(68912) := x"0062";
    tmp(68913) := x"0062";
    tmp(68914) := x"0062";
    tmp(68915) := x"0062";
    tmp(68916) := x"0062";
    tmp(68917) := x"0082";
    tmp(68918) := x"0062";
    tmp(68919) := x"0062";
    tmp(68920) := x"0041";
    tmp(68921) := x"0041";
    tmp(68922) := x"0041";
    tmp(68923) := x"0061";
    tmp(68924) := x"0062";
    tmp(68925) := x"0082";
    tmp(68926) := x"0062";
    tmp(68927) := x"0062";
    tmp(68928) := x"0062";
    tmp(68929) := x"0082";
    tmp(68930) := x"0062";
    tmp(68931) := x"0062";
    tmp(68932) := x"0061";
    tmp(68933) := x"0061";
    tmp(68934) := x"0062";
    tmp(68935) := x"0082";
    tmp(68936) := x"0082";
    tmp(68937) := x"0082";
    tmp(68938) := x"08a2";
    tmp(68939) := x"08a2";
    tmp(68940) := x"08a2";
    tmp(68941) := x"0081";
    tmp(68942) := x"0081";
    tmp(68943) := x"0040";
    tmp(68944) := x"0040";
    tmp(68945) := x"0040";
    tmp(68946) := x"0040";
    tmp(68947) := x"0040";
    tmp(68948) := x"0040";
    tmp(68949) := x"0040";
    tmp(68950) := x"0840";
    tmp(68951) := x"0840";
    tmp(68952) := x"0840";
    tmp(68953) := x"0020";
    tmp(68954) := x"0040";
    tmp(68955) := x"0840";
    tmp(68956) := x"0840";
    tmp(68957) := x"0840";
    tmp(68958) := x"0840";
    tmp(68959) := x"0820";
    tmp(68960) := x"0820";
    tmp(68961) := x"0820";
    tmp(68962) := x"0820";
    tmp(68963) := x"0820";
    tmp(68964) := x"0820";
    tmp(68965) := x"0820";
    tmp(68966) := x"0820";
    tmp(68967) := x"0820";
    tmp(68968) := x"0820";
    tmp(68969) := x"0820";
    tmp(68970) := x"1020";
    tmp(68971) := x"1000";
    tmp(68972) := x"1020";
    tmp(68973) := x"1820";
    tmp(68974) := x"1820";
    tmp(68975) := x"1020";
    tmp(68976) := x"0800";
    tmp(68977) := x"1000";
    tmp(68978) := x"1800";
    tmp(68979) := x"2000";
    tmp(68980) := x"2820";
    tmp(68981) := x"3000";
    tmp(68982) := x"3000";
    tmp(68983) := x"3800";
    tmp(68984) := x"3820";
    tmp(68985) := x"3000";
    tmp(68986) := x"3000";
    tmp(68987) := x"3000";
    tmp(68988) := x"3000";
    tmp(68989) := x"3820";
    tmp(68990) := x"3820";
    tmp(68991) := x"3020";
    tmp(68992) := x"2000";
    tmp(68993) := x"1000";
    tmp(68994) := x"0800";
    tmp(68995) := x"0800";
    tmp(68996) := x"1000";
    tmp(68997) := x"1800";
    tmp(68998) := x"2800";
    tmp(68999) := x"2800";
    tmp(69000) := x"3000";
    tmp(69001) := x"3000";
    tmp(69002) := x"2800";
    tmp(69003) := x"2000";
    tmp(69004) := x"1800";
    tmp(69005) := x"2000";
    tmp(69006) := x"2800";
    tmp(69007) := x"2800";
    tmp(69008) := x"2800";
    tmp(69009) := x"2800";
    tmp(69010) := x"3000";
    tmp(69011) := x"3800";
    tmp(69012) := x"3800";
    tmp(69013) := x"3800";
    tmp(69014) := x"3800";
    tmp(69015) := x"4000";
    tmp(69016) := x"4000";
    tmp(69017) := x"4000";
    tmp(69018) := x"4800";
    tmp(69019) := x"4000";
    tmp(69020) := x"4000";
    tmp(69021) := x"4000";
    tmp(69022) := x"4800";
    tmp(69023) := x"4000";
    tmp(69024) := x"3000";
    tmp(69025) := x"3000";
    tmp(69026) := x"5000";
    tmp(69027) := x"6020";
    tmp(69028) := x"5800";
    tmp(69029) := x"5020";
    tmp(69030) := x"4820";
    tmp(69031) := x"3081";
    tmp(69032) := x"3081";
    tmp(69033) := x"2061";
    tmp(69034) := x"20a1";
    tmp(69035) := x"20c2";
    tmp(69036) := x"20a2";
    tmp(69037) := x"18a2";
    tmp(69038) := x"18a2";
    tmp(69039) := x"18a2";
    tmp(69040) := x"18a2";
    tmp(69041) := x"18a1";
    tmp(69042) := x"18a1";
    tmp(69043) := x"18a1";
    tmp(69044) := x"1881";
    tmp(69045) := x"1081";
    tmp(69046) := x"1081";
    tmp(69047) := x"1061";
    tmp(69048) := x"1061";
    tmp(69049) := x"1061";
    tmp(69050) := x"1061";
    tmp(69051) := x"0840";
    tmp(69052) := x"0840";
    tmp(69053) := x"0840";
    tmp(69054) := x"0840";
    tmp(69055) := x"0840";
    tmp(69056) := x"0840";
    tmp(69057) := x"0840";
    tmp(69058) := x"0840";
    tmp(69059) := x"0820";
    tmp(69060) := x"0820";
    tmp(69061) := x"0820";
    tmp(69062) := x"0820";
    tmp(69063) := x"0820";
    tmp(69064) := x"0820";
    tmp(69065) := x"0840";
    tmp(69066) := x"0840";
    tmp(69067) := x"0841";
    tmp(69068) := x"0861";
    tmp(69069) := x"1081";
    tmp(69070) := x"1081";
    tmp(69071) := x"10a2";
    tmp(69072) := x"18c2";
    tmp(69073) := x"18e3";
    tmp(69074) := x"2104";
    tmp(69075) := x"2124";
    tmp(69076) := x"2144";
    tmp(69077) := x"2145";
    tmp(69078) := x"2945";
    tmp(69079) := x"2945";
    tmp(69080) := x"2966";
    tmp(69081) := x"3186";
    tmp(69082) := x"31a7";
    tmp(69083) := x"39c8";
    tmp(69084) := x"39e8";
    tmp(69085) := x"4209";
    tmp(69086) := x"4a2a";
    tmp(69087) := x"526b";
    tmp(69088) := x"5aad";
    tmp(69089) := x"5ace";
    tmp(69090) := x"6b4f";
    tmp(69091) := x"7370";
    tmp(69092) := x"7bb1";
    tmp(69093) := x"7bf2";
    tmp(69094) := x"83f3";
    tmp(69095) := x"83f3";
    tmp(69096) := x"83d3";
    tmp(69097) := x"7bb2";
    tmp(69098) := x"7bb2";
    tmp(69099) := x"7b92";
    tmp(69100) := x"7b92";
    tmp(69101) := x"7b72";
    tmp(69102) := x"7350";
    tmp(69103) := x"6b50";
    tmp(69104) := x"6b2f";
    tmp(69105) := x"6b4f";
    tmp(69106) := x"6b2f";
    tmp(69107) := x"6b0f";
    tmp(69108) := x"6b0f";
    tmp(69109) := x"62ee";
    tmp(69110) := x"5aee";
    tmp(69111) := x"5ace";
    tmp(69112) := x"5acd";
    tmp(69113) := x"5acd";
    tmp(69114) := x"52ad";
    tmp(69115) := x"528c";
    tmp(69116) := x"528b";
    tmp(69117) := x"4a6a";
    tmp(69118) := x"422a";
    tmp(69119) := x"4228";
    tmp(69120) := x"0000";
    tmp(69121) := x"0041";
    tmp(69122) := x"0041";
    tmp(69123) := x"0041";
    tmp(69124) := x"0041";
    tmp(69125) := x"0041";
    tmp(69126) := x"0041";
    tmp(69127) := x"0041";
    tmp(69128) := x"0041";
    tmp(69129) := x"0041";
    tmp(69130) := x"0041";
    tmp(69131) := x"0041";
    tmp(69132) := x"0041";
    tmp(69133) := x"0041";
    tmp(69134) := x"0041";
    tmp(69135) := x"0041";
    tmp(69136) := x"0041";
    tmp(69137) := x"0041";
    tmp(69138) := x"0041";
    tmp(69139) := x"0041";
    tmp(69140) := x"0041";
    tmp(69141) := x"0041";
    tmp(69142) := x"0041";
    tmp(69143) := x"0041";
    tmp(69144) := x"0041";
    tmp(69145) := x"0041";
    tmp(69146) := x"0041";
    tmp(69147) := x"0041";
    tmp(69148) := x"0041";
    tmp(69149) := x"0061";
    tmp(69150) := x"0062";
    tmp(69151) := x"0062";
    tmp(69152) := x"0062";
    tmp(69153) := x"0062";
    tmp(69154) := x"0062";
    tmp(69155) := x"0062";
    tmp(69156) := x"0062";
    tmp(69157) := x"0062";
    tmp(69158) := x"0062";
    tmp(69159) := x"0062";
    tmp(69160) := x"0062";
    tmp(69161) := x"0062";
    tmp(69162) := x"0062";
    tmp(69163) := x"0062";
    tmp(69164) := x"0062";
    tmp(69165) := x"0062";
    tmp(69166) := x"0061";
    tmp(69167) := x"0041";
    tmp(69168) := x"0041";
    tmp(69169) := x"0062";
    tmp(69170) := x"0062";
    tmp(69171) := x"0062";
    tmp(69172) := x"0062";
    tmp(69173) := x"0082";
    tmp(69174) := x"0082";
    tmp(69175) := x"00a2";
    tmp(69176) := x"00a2";
    tmp(69177) := x"08a2";
    tmp(69178) := x"0082";
    tmp(69179) := x"0081";
    tmp(69180) := x"0061";
    tmp(69181) := x"0061";
    tmp(69182) := x"0061";
    tmp(69183) := x"0040";
    tmp(69184) := x"0040";
    tmp(69185) := x"0040";
    tmp(69186) := x"0040";
    tmp(69187) := x"0040";
    tmp(69188) := x"0040";
    tmp(69189) := x"0040";
    tmp(69190) := x"0040";
    tmp(69191) := x"0840";
    tmp(69192) := x"0820";
    tmp(69193) := x"0820";
    tmp(69194) := x"0820";
    tmp(69195) := x"0820";
    tmp(69196) := x"0820";
    tmp(69197) := x"0820";
    tmp(69198) := x"0820";
    tmp(69199) := x"0820";
    tmp(69200) := x"0820";
    tmp(69201) := x"0820";
    tmp(69202) := x"0820";
    tmp(69203) := x"0820";
    tmp(69204) := x"1020";
    tmp(69205) := x"1020";
    tmp(69206) := x"1020";
    tmp(69207) := x"0820";
    tmp(69208) := x"0820";
    tmp(69209) := x"1000";
    tmp(69210) := x"1820";
    tmp(69211) := x"1820";
    tmp(69212) := x"2020";
    tmp(69213) := x"2020";
    tmp(69214) := x"1820";
    tmp(69215) := x"1000";
    tmp(69216) := x"1000";
    tmp(69217) := x"1800";
    tmp(69218) := x"2000";
    tmp(69219) := x"2820";
    tmp(69220) := x"3020";
    tmp(69221) := x"3020";
    tmp(69222) := x"3000";
    tmp(69223) := x"3000";
    tmp(69224) := x"3800";
    tmp(69225) := x"3000";
    tmp(69226) := x"3000";
    tmp(69227) := x"3800";
    tmp(69228) := x"3820";
    tmp(69229) := x"4020";
    tmp(69230) := x"4020";
    tmp(69231) := x"3020";
    tmp(69232) := x"2000";
    tmp(69233) := x"1000";
    tmp(69234) := x"1000";
    tmp(69235) := x"1000";
    tmp(69236) := x"1000";
    tmp(69237) := x"1000";
    tmp(69238) := x"1800";
    tmp(69239) := x"2800";
    tmp(69240) := x"3000";
    tmp(69241) := x"2800";
    tmp(69242) := x"2000";
    tmp(69243) := x"1800";
    tmp(69244) := x"2000";
    tmp(69245) := x"3000";
    tmp(69246) := x"3000";
    tmp(69247) := x"2800";
    tmp(69248) := x"2800";
    tmp(69249) := x"3000";
    tmp(69250) := x"3800";
    tmp(69251) := x"3800";
    tmp(69252) := x"4800";
    tmp(69253) := x"3800";
    tmp(69254) := x"3800";
    tmp(69255) := x"3800";
    tmp(69256) := x"3800";
    tmp(69257) := x"4000";
    tmp(69258) := x"4000";
    tmp(69259) := x"4000";
    tmp(69260) := x"4000";
    tmp(69261) := x"4000";
    tmp(69262) := x"4000";
    tmp(69263) := x"3800";
    tmp(69264) := x"2800";
    tmp(69265) := x"4000";
    tmp(69266) := x"6820";
    tmp(69267) := x"6020";
    tmp(69268) := x"4000";
    tmp(69269) := x"4820";
    tmp(69270) := x"3061";
    tmp(69271) := x"20a1";
    tmp(69272) := x"2081";
    tmp(69273) := x"18a1";
    tmp(69274) := x"18a1";
    tmp(69275) := x"18a1";
    tmp(69276) := x"18a2";
    tmp(69277) := x"18a2";
    tmp(69278) := x"18a1";
    tmp(69279) := x"18a1";
    tmp(69280) := x"18a1";
    tmp(69281) := x"18a1";
    tmp(69282) := x"18a1";
    tmp(69283) := x"1881";
    tmp(69284) := x"1081";
    tmp(69285) := x"1081";
    tmp(69286) := x"1061";
    tmp(69287) := x"1061";
    tmp(69288) := x"1061";
    tmp(69289) := x"1061";
    tmp(69290) := x"1061";
    tmp(69291) := x"0840";
    tmp(69292) := x"0840";
    tmp(69293) := x"0840";
    tmp(69294) := x"0840";
    tmp(69295) := x"0840";
    tmp(69296) := x"0840";
    tmp(69297) := x"0840";
    tmp(69298) := x"0820";
    tmp(69299) := x"0820";
    tmp(69300) := x"0820";
    tmp(69301) := x"0820";
    tmp(69302) := x"0820";
    tmp(69303) := x"0820";
    tmp(69304) := x"0820";
    tmp(69305) := x"0840";
    tmp(69306) := x"0840";
    tmp(69307) := x"0841";
    tmp(69308) := x"0841";
    tmp(69309) := x"0861";
    tmp(69310) := x"1081";
    tmp(69311) := x"1081";
    tmp(69312) := x"10a2";
    tmp(69313) := x"18c2";
    tmp(69314) := x"18c3";
    tmp(69315) := x"18e3";
    tmp(69316) := x"1903";
    tmp(69317) := x"2103";
    tmp(69318) := x"2104";
    tmp(69319) := x"2124";
    tmp(69320) := x"2925";
    tmp(69321) := x"2965";
    tmp(69322) := x"3186";
    tmp(69323) := x"3186";
    tmp(69324) := x"31a7";
    tmp(69325) := x"39c8";
    tmp(69326) := x"39e9";
    tmp(69327) := x"422a";
    tmp(69328) := x"4a4a";
    tmp(69329) := x"52ad";
    tmp(69330) := x"5acd";
    tmp(69331) := x"630e";
    tmp(69332) := x"6b4f";
    tmp(69333) := x"7371";
    tmp(69334) := x"7371";
    tmp(69335) := x"7391";
    tmp(69336) := x"7b91";
    tmp(69337) := x"7371";
    tmp(69338) := x"7371";
    tmp(69339) := x"7370";
    tmp(69340) := x"7351";
    tmp(69341) := x"6b30";
    tmp(69342) := x"6b30";
    tmp(69343) := x"6b0f";
    tmp(69344) := x"6b2f";
    tmp(69345) := x"630f";
    tmp(69346) := x"630f";
    tmp(69347) := x"630f";
    tmp(69348) := x"62ee";
    tmp(69349) := x"5aee";
    tmp(69350) := x"5ace";
    tmp(69351) := x"5aad";
    tmp(69352) := x"528d";
    tmp(69353) := x"528d";
    tmp(69354) := x"528c";
    tmp(69355) := x"526c";
    tmp(69356) := x"526b";
    tmp(69357) := x"4a4a";
    tmp(69358) := x"4229";
    tmp(69359) := x"39e8";
    tmp(69360) := x"0000";
    tmp(69361) := x"0041";
    tmp(69362) := x"0041";
    tmp(69363) := x"0041";
    tmp(69364) := x"0041";
    tmp(69365) := x"0041";
    tmp(69366) := x"0041";
    tmp(69367) := x"0041";
    tmp(69368) := x"0041";
    tmp(69369) := x"0041";
    tmp(69370) := x"0041";
    tmp(69371) := x"0041";
    tmp(69372) := x"0041";
    tmp(69373) := x"0041";
    tmp(69374) := x"0041";
    tmp(69375) := x"0041";
    tmp(69376) := x"0041";
    tmp(69377) := x"0041";
    tmp(69378) := x"0041";
    tmp(69379) := x"0041";
    tmp(69380) := x"0061";
    tmp(69381) := x"0061";
    tmp(69382) := x"0061";
    tmp(69383) := x"0041";
    tmp(69384) := x"0041";
    tmp(69385) := x"0041";
    tmp(69386) := x"0041";
    tmp(69387) := x"0041";
    tmp(69388) := x"0041";
    tmp(69389) := x"0041";
    tmp(69390) := x"0061";
    tmp(69391) := x"0061";
    tmp(69392) := x"0062";
    tmp(69393) := x"0062";
    tmp(69394) := x"0062";
    tmp(69395) := x"0062";
    tmp(69396) := x"0062";
    tmp(69397) := x"0062";
    tmp(69398) := x"0062";
    tmp(69399) := x"0062";
    tmp(69400) := x"0061";
    tmp(69401) := x"0061";
    tmp(69402) := x"0062";
    tmp(69403) := x"0041";
    tmp(69404) := x"0041";
    tmp(69405) := x"0041";
    tmp(69406) := x"0041";
    tmp(69407) := x"0061";
    tmp(69408) := x"0061";
    tmp(69409) := x"0082";
    tmp(69410) := x"0082";
    tmp(69411) := x"00a2";
    tmp(69412) := x"00a2";
    tmp(69413) := x"00a2";
    tmp(69414) := x"00a2";
    tmp(69415) := x"0082";
    tmp(69416) := x"0081";
    tmp(69417) := x"0081";
    tmp(69418) := x"0061";
    tmp(69419) := x"0061";
    tmp(69420) := x"0061";
    tmp(69421) := x"0061";
    tmp(69422) := x"0061";
    tmp(69423) := x"0060";
    tmp(69424) := x"0040";
    tmp(69425) := x"0040";
    tmp(69426) := x"0040";
    tmp(69427) := x"0040";
    tmp(69428) := x"0040";
    tmp(69429) := x"0020";
    tmp(69430) := x"0020";
    tmp(69431) := x"0020";
    tmp(69432) := x"0020";
    tmp(69433) := x"0020";
    tmp(69434) := x"0820";
    tmp(69435) := x"0820";
    tmp(69436) := x"0800";
    tmp(69437) := x"0800";
    tmp(69438) := x"1000";
    tmp(69439) := x"1000";
    tmp(69440) := x"1000";
    tmp(69441) := x"1000";
    tmp(69442) := x"1000";
    tmp(69443) := x"1000";
    tmp(69444) := x"1000";
    tmp(69445) := x"1820";
    tmp(69446) := x"1020";
    tmp(69447) := x"1020";
    tmp(69448) := x"1020";
    tmp(69449) := x"1800";
    tmp(69450) := x"2020";
    tmp(69451) := x"2820";
    tmp(69452) := x"2820";
    tmp(69453) := x"2820";
    tmp(69454) := x"2020";
    tmp(69455) := x"1000";
    tmp(69456) := x"1800";
    tmp(69457) := x"2000";
    tmp(69458) := x"2800";
    tmp(69459) := x"3000";
    tmp(69460) := x"3020";
    tmp(69461) := x"3020";
    tmp(69462) := x"3000";
    tmp(69463) := x"3000";
    tmp(69464) := x"3800";
    tmp(69465) := x"3000";
    tmp(69466) := x"3000";
    tmp(69467) := x"3800";
    tmp(69468) := x"4020";
    tmp(69469) := x"4820";
    tmp(69470) := x"5020";
    tmp(69471) := x"3820";
    tmp(69472) := x"2000";
    tmp(69473) := x"1800";
    tmp(69474) := x"1800";
    tmp(69475) := x"2000";
    tmp(69476) := x"1800";
    tmp(69477) := x"1000";
    tmp(69478) := x"1800";
    tmp(69479) := x"2800";
    tmp(69480) := x"2800";
    tmp(69481) := x"2000";
    tmp(69482) := x"1800";
    tmp(69483) := x"2000";
    tmp(69484) := x"2800";
    tmp(69485) := x"3000";
    tmp(69486) := x"3000";
    tmp(69487) := x"3000";
    tmp(69488) := x"3000";
    tmp(69489) := x"3000";
    tmp(69490) := x"3800";
    tmp(69491) := x"4800";
    tmp(69492) := x"4000";
    tmp(69493) := x"3800";
    tmp(69494) := x"3000";
    tmp(69495) := x"3000";
    tmp(69496) := x"3800";
    tmp(69497) := x"3800";
    tmp(69498) := x"3800";
    tmp(69499) := x"3800";
    tmp(69500) := x"4000";
    tmp(69501) := x"4000";
    tmp(69502) := x"3000";
    tmp(69503) := x"2000";
    tmp(69504) := x"2800";
    tmp(69505) := x"5020";
    tmp(69506) := x"5820";
    tmp(69507) := x"5020";
    tmp(69508) := x"5020";
    tmp(69509) := x"4041";
    tmp(69510) := x"20a1";
    tmp(69511) := x"18a1";
    tmp(69512) := x"18a1";
    tmp(69513) := x"18a1";
    tmp(69514) := x"18a1";
    tmp(69515) := x"18a1";
    tmp(69516) := x"18a1";
    tmp(69517) := x"18a1";
    tmp(69518) := x"18a1";
    tmp(69519) := x"18a1";
    tmp(69520) := x"18a1";
    tmp(69521) := x"18a1";
    tmp(69522) := x"18a1";
    tmp(69523) := x"1881";
    tmp(69524) := x"1081";
    tmp(69525) := x"1081";
    tmp(69526) := x"1061";
    tmp(69527) := x"1061";
    tmp(69528) := x"1061";
    tmp(69529) := x"1061";
    tmp(69530) := x"1061";
    tmp(69531) := x"0840";
    tmp(69532) := x"0840";
    tmp(69533) := x"0840";
    tmp(69534) := x"0840";
    tmp(69535) := x"0840";
    tmp(69536) := x"0840";
    tmp(69537) := x"0820";
    tmp(69538) := x"0820";
    tmp(69539) := x"0820";
    tmp(69540) := x"0820";
    tmp(69541) := x"0820";
    tmp(69542) := x"0820";
    tmp(69543) := x"0820";
    tmp(69544) := x"0820";
    tmp(69545) := x"0820";
    tmp(69546) := x"0820";
    tmp(69547) := x"0840";
    tmp(69548) := x"0841";
    tmp(69549) := x"0841";
    tmp(69550) := x"0861";
    tmp(69551) := x"1061";
    tmp(69552) := x"1081";
    tmp(69553) := x"1081";
    tmp(69554) := x"10a2";
    tmp(69555) := x"10a2";
    tmp(69556) := x"18c2";
    tmp(69557) := x"18c3";
    tmp(69558) := x"18e3";
    tmp(69559) := x"18e3";
    tmp(69560) := x"2104";
    tmp(69561) := x"2124";
    tmp(69562) := x"2945";
    tmp(69563) := x"2965";
    tmp(69564) := x"2966";
    tmp(69565) := x"3186";
    tmp(69566) := x"39a7";
    tmp(69567) := x"39e8";
    tmp(69568) := x"4209";
    tmp(69569) := x"4a6b";
    tmp(69570) := x"528b";
    tmp(69571) := x"5aed";
    tmp(69572) := x"630e";
    tmp(69573) := x"630e";
    tmp(69574) := x"6b0e";
    tmp(69575) := x"6b4f";
    tmp(69576) := x"6b2f";
    tmp(69577) := x"6b50";
    tmp(69578) := x"6b4f";
    tmp(69579) := x"6b2f";
    tmp(69580) := x"6b2f";
    tmp(69581) := x"6b0f";
    tmp(69582) := x"6b0f";
    tmp(69583) := x"62cf";
    tmp(69584) := x"62ef";
    tmp(69585) := x"5ace";
    tmp(69586) := x"5ace";
    tmp(69587) := x"62ce";
    tmp(69588) := x"5acd";
    tmp(69589) := x"5acd";
    tmp(69590) := x"5acd";
    tmp(69591) := x"5aad";
    tmp(69592) := x"526c";
    tmp(69593) := x"526c";
    tmp(69594) := x"4a4b";
    tmp(69595) := x"4a4b";
    tmp(69596) := x"4a4b";
    tmp(69597) := x"422a";
    tmp(69598) := x"3a08";
    tmp(69599) := x"39e8";
    tmp(69600) := x"0000";
    tmp(69601) := x"0041";
    tmp(69602) := x"0041";
    tmp(69603) := x"0041";
    tmp(69604) := x"0041";
    tmp(69605) := x"0041";
    tmp(69606) := x"0041";
    tmp(69607) := x"0041";
    tmp(69608) := x"0041";
    tmp(69609) := x"0041";
    tmp(69610) := x"0041";
    tmp(69611) := x"0041";
    tmp(69612) := x"0041";
    tmp(69613) := x"0041";
    tmp(69614) := x"0041";
    tmp(69615) := x"0041";
    tmp(69616) := x"0041";
    tmp(69617) := x"0041";
    tmp(69618) := x"0041";
    tmp(69619) := x"0041";
    tmp(69620) := x"0041";
    tmp(69621) := x"0041";
    tmp(69622) := x"0061";
    tmp(69623) := x"0061";
    tmp(69624) := x"0061";
    tmp(69625) := x"0041";
    tmp(69626) := x"0061";
    tmp(69627) := x"0041";
    tmp(69628) := x"0041";
    tmp(69629) := x"0041";
    tmp(69630) := x"0041";
    tmp(69631) := x"0041";
    tmp(69632) := x"0041";
    tmp(69633) := x"0041";
    tmp(69634) := x"0061";
    tmp(69635) := x"0061";
    tmp(69636) := x"0061";
    tmp(69637) := x"0062";
    tmp(69638) := x"0062";
    tmp(69639) := x"0062";
    tmp(69640) := x"0062";
    tmp(69641) := x"0062";
    tmp(69642) := x"0061";
    tmp(69643) := x"0041";
    tmp(69644) := x"0041";
    tmp(69645) := x"0041";
    tmp(69646) := x"0061";
    tmp(69647) := x"0061";
    tmp(69648) := x"0061";
    tmp(69649) := x"0082";
    tmp(69650) := x"0082";
    tmp(69651) := x"0082";
    tmp(69652) := x"0082";
    tmp(69653) := x"0082";
    tmp(69654) := x"0081";
    tmp(69655) := x"0061";
    tmp(69656) := x"0061";
    tmp(69657) := x"0061";
    tmp(69658) := x"0061";
    tmp(69659) := x"0061";
    tmp(69660) := x"0061";
    tmp(69661) := x"0061";
    tmp(69662) := x"0061";
    tmp(69663) := x"0060";
    tmp(69664) := x"0060";
    tmp(69665) := x"0060";
    tmp(69666) := x"0040";
    tmp(69667) := x"0840";
    tmp(69668) := x"0040";
    tmp(69669) := x"0020";
    tmp(69670) := x"0020";
    tmp(69671) := x"0020";
    tmp(69672) := x"0020";
    tmp(69673) := x"0020";
    tmp(69674) := x"0820";
    tmp(69675) := x"0820";
    tmp(69676) := x"1000";
    tmp(69677) := x"1000";
    tmp(69678) := x"1800";
    tmp(69679) := x"1800";
    tmp(69680) := x"1800";
    tmp(69681) := x"1800";
    tmp(69682) := x"1800";
    tmp(69683) := x"1800";
    tmp(69684) := x"1800";
    tmp(69685) := x"1800";
    tmp(69686) := x"1000";
    tmp(69687) := x"1000";
    tmp(69688) := x"1000";
    tmp(69689) := x"1800";
    tmp(69690) := x"2000";
    tmp(69691) := x"2800";
    tmp(69692) := x"2800";
    tmp(69693) := x"3020";
    tmp(69694) := x"2820";
    tmp(69695) := x"2000";
    tmp(69696) := x"2000";
    tmp(69697) := x"2800";
    tmp(69698) := x"2800";
    tmp(69699) := x"3000";
    tmp(69700) := x"3020";
    tmp(69701) := x"3820";
    tmp(69702) := x"3820";
    tmp(69703) := x"2800";
    tmp(69704) := x"3000";
    tmp(69705) := x"3000";
    tmp(69706) := x"4020";
    tmp(69707) := x"4020";
    tmp(69708) := x"4820";
    tmp(69709) := x"5020";
    tmp(69710) := x"5020";
    tmp(69711) := x"3820";
    tmp(69712) := x"3000";
    tmp(69713) := x"3000";
    tmp(69714) := x"3000";
    tmp(69715) := x"2000";
    tmp(69716) := x"1000";
    tmp(69717) := x"2020";
    tmp(69718) := x"2000";
    tmp(69719) := x"2800";
    tmp(69720) := x"1800";
    tmp(69721) := x"1800";
    tmp(69722) := x"2000";
    tmp(69723) := x"2000";
    tmp(69724) := x"3000";
    tmp(69725) := x"3800";
    tmp(69726) := x"3800";
    tmp(69727) := x"3800";
    tmp(69728) := x"3800";
    tmp(69729) := x"3800";
    tmp(69730) := x"4000";
    tmp(69731) := x"4000";
    tmp(69732) := x"4820";
    tmp(69733) := x"3000";
    tmp(69734) := x"3820";
    tmp(69735) := x"3020";
    tmp(69736) := x"2800";
    tmp(69737) := x"2800";
    tmp(69738) := x"3000";
    tmp(69739) := x"3000";
    tmp(69740) := x"3800";
    tmp(69741) := x"3800";
    tmp(69742) := x"2000";
    tmp(69743) := x"1800";
    tmp(69744) := x"3820";
    tmp(69745) := x"6020";
    tmp(69746) := x"5820";
    tmp(69747) := x"4820";
    tmp(69748) := x"4861";
    tmp(69749) := x"2881";
    tmp(69750) := x"18a1";
    tmp(69751) := x"18a1";
    tmp(69752) := x"18a1";
    tmp(69753) := x"18a1";
    tmp(69754) := x"18a1";
    tmp(69755) := x"18a1";
    tmp(69756) := x"18a1";
    tmp(69757) := x"18a1";
    tmp(69758) := x"18a1";
    tmp(69759) := x"18a1";
    tmp(69760) := x"18a1";
    tmp(69761) := x"18a1";
    tmp(69762) := x"1081";
    tmp(69763) := x"1081";
    tmp(69764) := x"1081";
    tmp(69765) := x"1081";
    tmp(69766) := x"1061";
    tmp(69767) := x"1061";
    tmp(69768) := x"1061";
    tmp(69769) := x"1061";
    tmp(69770) := x"0861";
    tmp(69771) := x"0840";
    tmp(69772) := x"0840";
    tmp(69773) := x"0840";
    tmp(69774) := x"0840";
    tmp(69775) := x"0840";
    tmp(69776) := x"0840";
    tmp(69777) := x"0840";
    tmp(69778) := x"0820";
    tmp(69779) := x"0820";
    tmp(69780) := x"0820";
    tmp(69781) := x"0820";
    tmp(69782) := x"0820";
    tmp(69783) := x"0820";
    tmp(69784) := x"0820";
    tmp(69785) := x"0820";
    tmp(69786) := x"0820";
    tmp(69787) := x"0820";
    tmp(69788) := x"0840";
    tmp(69789) := x"0841";
    tmp(69790) := x"0841";
    tmp(69791) := x"0861";
    tmp(69792) := x"0861";
    tmp(69793) := x"1061";
    tmp(69794) := x"1081";
    tmp(69795) := x"1081";
    tmp(69796) := x"10a2";
    tmp(69797) := x"10a2";
    tmp(69798) := x"18c2";
    tmp(69799) := x"18c2";
    tmp(69800) := x"18c3";
    tmp(69801) := x"18e3";
    tmp(69802) := x"2104";
    tmp(69803) := x"2124";
    tmp(69804) := x"2124";
    tmp(69805) := x"2945";
    tmp(69806) := x"3186";
    tmp(69807) := x"31a7";
    tmp(69808) := x"31a7";
    tmp(69809) := x"3a08";
    tmp(69810) := x"4a49";
    tmp(69811) := x"526a";
    tmp(69812) := x"5acb";
    tmp(69813) := x"5aac";
    tmp(69814) := x"62cd";
    tmp(69815) := x"62ee";
    tmp(69816) := x"5ace";
    tmp(69817) := x"62ee";
    tmp(69818) := x"62ee";
    tmp(69819) := x"62ce";
    tmp(69820) := x"62ce";
    tmp(69821) := x"62ef";
    tmp(69822) := x"62cf";
    tmp(69823) := x"5aae";
    tmp(69824) := x"5acd";
    tmp(69825) := x"5aad";
    tmp(69826) := x"5acd";
    tmp(69827) := x"5aad";
    tmp(69828) := x"5aad";
    tmp(69829) := x"5aae";
    tmp(69830) := x"52ad";
    tmp(69831) := x"528d";
    tmp(69832) := x"526c";
    tmp(69833) := x"4a4b";
    tmp(69834) := x"4a4b";
    tmp(69835) := x"424a";
    tmp(69836) := x"422a";
    tmp(69837) := x"4209";
    tmp(69838) := x"39c8";
    tmp(69839) := x"39c7";
    tmp(69840) := x"0000";
    tmp(69841) := x"0041";
    tmp(69842) := x"0041";
    tmp(69843) := x"0041";
    tmp(69844) := x"0041";
    tmp(69845) := x"0041";
    tmp(69846) := x"0041";
    tmp(69847) := x"0041";
    tmp(69848) := x"0041";
    tmp(69849) := x"0041";
    tmp(69850) := x"0041";
    tmp(69851) := x"0041";
    tmp(69852) := x"0041";
    tmp(69853) := x"0041";
    tmp(69854) := x"0041";
    tmp(69855) := x"0041";
    tmp(69856) := x"0041";
    tmp(69857) := x"0041";
    tmp(69858) := x"0041";
    tmp(69859) := x"0041";
    tmp(69860) := x"0041";
    tmp(69861) := x"0041";
    tmp(69862) := x"0061";
    tmp(69863) := x"0061";
    tmp(69864) := x"0061";
    tmp(69865) := x"0041";
    tmp(69866) := x"0061";
    tmp(69867) := x"0061";
    tmp(69868) := x"0061";
    tmp(69869) := x"0061";
    tmp(69870) := x"0061";
    tmp(69871) := x"0041";
    tmp(69872) := x"0041";
    tmp(69873) := x"0041";
    tmp(69874) := x"0041";
    tmp(69875) := x"0041";
    tmp(69876) := x"0041";
    tmp(69877) := x"0041";
    tmp(69878) := x"0062";
    tmp(69879) := x"0062";
    tmp(69880) := x"0062";
    tmp(69881) := x"0062";
    tmp(69882) := x"0041";
    tmp(69883) := x"0041";
    tmp(69884) := x"0041";
    tmp(69885) := x"0041";
    tmp(69886) := x"0061";
    tmp(69887) := x"0061";
    tmp(69888) := x"0061";
    tmp(69889) := x"0061";
    tmp(69890) := x"0061";
    tmp(69891) := x"0061";
    tmp(69892) := x"0061";
    tmp(69893) := x"0061";
    tmp(69894) := x"0061";
    tmp(69895) := x"0061";
    tmp(69896) := x"0061";
    tmp(69897) := x"0061";
    tmp(69898) := x"0060";
    tmp(69899) := x"0060";
    tmp(69900) := x"0061";
    tmp(69901) := x"0061";
    tmp(69902) := x"0060";
    tmp(69903) := x"0060";
    tmp(69904) := x"0060";
    tmp(69905) := x"0060";
    tmp(69906) := x"0860";
    tmp(69907) := x"0860";
    tmp(69908) := x"0840";
    tmp(69909) := x"0840";
    tmp(69910) := x"0820";
    tmp(69911) := x"0820";
    tmp(69912) := x"0020";
    tmp(69913) := x"0020";
    tmp(69914) := x"0000";
    tmp(69915) := x"0800";
    tmp(69916) := x"0800";
    tmp(69917) := x"1000";
    tmp(69918) := x"1800";
    tmp(69919) := x"2000";
    tmp(69920) := x"2000";
    tmp(69921) := x"2000";
    tmp(69922) := x"1800";
    tmp(69923) := x"1800";
    tmp(69924) := x"1800";
    tmp(69925) := x"1800";
    tmp(69926) := x"1000";
    tmp(69927) := x"1000";
    tmp(69928) := x"1800";
    tmp(69929) := x"1800";
    tmp(69930) := x"2000";
    tmp(69931) := x"2800";
    tmp(69932) := x"2820";
    tmp(69933) := x"2820";
    tmp(69934) := x"2820";
    tmp(69935) := x"2020";
    tmp(69936) := x"2000";
    tmp(69937) := x"2800";
    tmp(69938) := x"3000";
    tmp(69939) := x"3000";
    tmp(69940) := x"3820";
    tmp(69941) := x"3820";
    tmp(69942) := x"3020";
    tmp(69943) := x"2800";
    tmp(69944) := x"3000";
    tmp(69945) := x"3000";
    tmp(69946) := x"4020";
    tmp(69947) := x"3820";
    tmp(69948) := x"4020";
    tmp(69949) := x"4020";
    tmp(69950) := x"4020";
    tmp(69951) := x"3800";
    tmp(69952) := x"3800";
    tmp(69953) := x"4820";
    tmp(69954) := x"4020";
    tmp(69955) := x"1800";
    tmp(69956) := x"0800";
    tmp(69957) := x"2820";
    tmp(69958) := x"2800";
    tmp(69959) := x"2800";
    tmp(69960) := x"1800";
    tmp(69961) := x"1800";
    tmp(69962) := x"2000";
    tmp(69963) := x"2800";
    tmp(69964) := x"3000";
    tmp(69965) := x"3800";
    tmp(69966) := x"4000";
    tmp(69967) := x"3800";
    tmp(69968) := x"3800";
    tmp(69969) := x"3000";
    tmp(69970) := x"2800";
    tmp(69971) := x"4020";
    tmp(69972) := x"3020";
    tmp(69973) := x"2800";
    tmp(69974) := x"3020";
    tmp(69975) := x"1800";
    tmp(69976) := x"1800";
    tmp(69977) := x"2800";
    tmp(69978) := x"3820";
    tmp(69979) := x"3000";
    tmp(69980) := x"3000";
    tmp(69981) := x"2800";
    tmp(69982) := x"1800";
    tmp(69983) := x"1800";
    tmp(69984) := x"4820";
    tmp(69985) := x"5840";
    tmp(69986) := x"4841";
    tmp(69987) := x"3881";
    tmp(69988) := x"2881";
    tmp(69989) := x"18a1";
    tmp(69990) := x"18a1";
    tmp(69991) := x"18a1";
    tmp(69992) := x"18a1";
    tmp(69993) := x"18a1";
    tmp(69994) := x"18a1";
    tmp(69995) := x"1881";
    tmp(69996) := x"1881";
    tmp(69997) := x"1081";
    tmp(69998) := x"1081";
    tmp(69999) := x"1081";
    tmp(70000) := x"1081";
    tmp(70001) := x"1081";
    tmp(70002) := x"1081";
    tmp(70003) := x"1081";
    tmp(70004) := x"1081";
    tmp(70005) := x"1061";
    tmp(70006) := x"1061";
    tmp(70007) := x"1061";
    tmp(70008) := x"1061";
    tmp(70009) := x"1061";
    tmp(70010) := x"0840";
    tmp(70011) := x"0840";
    tmp(70012) := x"0840";
    tmp(70013) := x"0840";
    tmp(70014) := x"0840";
    tmp(70015) := x"0840";
    tmp(70016) := x"0840";
    tmp(70017) := x"0840";
    tmp(70018) := x"0820";
    tmp(70019) := x"0820";
    tmp(70020) := x"0820";
    tmp(70021) := x"0820";
    tmp(70022) := x"0820";
    tmp(70023) := x"0820";
    tmp(70024) := x"0820";
    tmp(70025) := x"0820";
    tmp(70026) := x"0820";
    tmp(70027) := x"0820";
    tmp(70028) := x"0820";
    tmp(70029) := x"0840";
    tmp(70030) := x"0840";
    tmp(70031) := x"0841";
    tmp(70032) := x"0841";
    tmp(70033) := x"0841";
    tmp(70034) := x"0861";
    tmp(70035) := x"0861";
    tmp(70036) := x"1061";
    tmp(70037) := x"1081";
    tmp(70038) := x"10a1";
    tmp(70039) := x"10a2";
    tmp(70040) := x"10a2";
    tmp(70041) := x"18c2";
    tmp(70042) := x"18e3";
    tmp(70043) := x"18e3";
    tmp(70044) := x"18e3";
    tmp(70045) := x"2104";
    tmp(70046) := x"2944";
    tmp(70047) := x"2965";
    tmp(70048) := x"3186";
    tmp(70049) := x"31a6";
    tmp(70050) := x"39e7";
    tmp(70051) := x"4208";
    tmp(70052) := x"4a49";
    tmp(70053) := x"526a";
    tmp(70054) := x"528c";
    tmp(70055) := x"528c";
    tmp(70056) := x"528c";
    tmp(70057) := x"5acd";
    tmp(70058) := x"5acd";
    tmp(70059) := x"5aad";
    tmp(70060) := x"5aad";
    tmp(70061) := x"5acd";
    tmp(70062) := x"5aad";
    tmp(70063) := x"5aad";
    tmp(70064) := x"5aad";
    tmp(70065) := x"526c";
    tmp(70066) := x"528c";
    tmp(70067) := x"528c";
    tmp(70068) := x"528d";
    tmp(70069) := x"526c";
    tmp(70070) := x"528d";
    tmp(70071) := x"526c";
    tmp(70072) := x"4a4b";
    tmp(70073) := x"4a4a";
    tmp(70074) := x"422a";
    tmp(70075) := x"4229";
    tmp(70076) := x"3a09";
    tmp(70077) := x"39e8";
    tmp(70078) := x"31a7";
    tmp(70079) := x"3186";
    tmp(70080) := x"0000";
    tmp(70081) := x"0041";
    tmp(70082) := x"0041";
    tmp(70083) := x"0041";
    tmp(70084) := x"0041";
    tmp(70085) := x"0041";
    tmp(70086) := x"0041";
    tmp(70087) := x"0041";
    tmp(70088) := x"0041";
    tmp(70089) := x"0041";
    tmp(70090) := x"0041";
    tmp(70091) := x"0041";
    tmp(70092) := x"0041";
    tmp(70093) := x"0041";
    tmp(70094) := x"0041";
    tmp(70095) := x"0041";
    tmp(70096) := x"0041";
    tmp(70097) := x"0041";
    tmp(70098) := x"0041";
    tmp(70099) := x"0041";
    tmp(70100) := x"0041";
    tmp(70101) := x"0041";
    tmp(70102) := x"0061";
    tmp(70103) := x"0061";
    tmp(70104) := x"0041";
    tmp(70105) := x"0061";
    tmp(70106) := x"0041";
    tmp(70107) := x"0061";
    tmp(70108) := x"0061";
    tmp(70109) := x"0061";
    tmp(70110) := x"0061";
    tmp(70111) := x"0062";
    tmp(70112) := x"0061";
    tmp(70113) := x"0041";
    tmp(70114) := x"0041";
    tmp(70115) := x"0041";
    tmp(70116) := x"0061";
    tmp(70117) := x"0062";
    tmp(70118) := x"0062";
    tmp(70119) := x"0062";
    tmp(70120) := x"0062";
    tmp(70121) := x"0062";
    tmp(70122) := x"0041";
    tmp(70123) := x"0041";
    tmp(70124) := x"0041";
    tmp(70125) := x"0041";
    tmp(70126) := x"0061";
    tmp(70127) := x"0041";
    tmp(70128) := x"0041";
    tmp(70129) := x"0061";
    tmp(70130) := x"0061";
    tmp(70131) := x"0061";
    tmp(70132) := x"0061";
    tmp(70133) := x"0061";
    tmp(70134) := x"0061";
    tmp(70135) := x"0061";
    tmp(70136) := x"0061";
    tmp(70137) := x"0061";
    tmp(70138) := x"0060";
    tmp(70139) := x"0060";
    tmp(70140) := x"0061";
    tmp(70141) := x"0061";
    tmp(70142) := x"0081";
    tmp(70143) := x"0060";
    tmp(70144) := x"0060";
    tmp(70145) := x"0880";
    tmp(70146) := x"0880";
    tmp(70147) := x"0881";
    tmp(70148) := x"0840";
    tmp(70149) := x"0840";
    tmp(70150) := x"0820";
    tmp(70151) := x"0820";
    tmp(70152) := x"0820";
    tmp(70153) := x"0820";
    tmp(70154) := x"0020";
    tmp(70155) := x"0000";
    tmp(70156) := x"0000";
    tmp(70157) := x"0800";
    tmp(70158) := x"1000";
    tmp(70159) := x"1800";
    tmp(70160) := x"2000";
    tmp(70161) := x"2000";
    tmp(70162) := x"2000";
    tmp(70163) := x"2000";
    tmp(70164) := x"1800";
    tmp(70165) := x"1800";
    tmp(70166) := x"1000";
    tmp(70167) := x"1000";
    tmp(70168) := x"1800";
    tmp(70169) := x"2000";
    tmp(70170) := x"2000";
    tmp(70171) := x"2000";
    tmp(70172) := x"2000";
    tmp(70173) := x"2000";
    tmp(70174) := x"2020";
    tmp(70175) := x"2000";
    tmp(70176) := x"2000";
    tmp(70177) := x"2800";
    tmp(70178) := x"3000";
    tmp(70179) := x"3800";
    tmp(70180) := x"3820";
    tmp(70181) := x"3820";
    tmp(70182) := x"2800";
    tmp(70183) := x"2800";
    tmp(70184) := x"2800";
    tmp(70185) := x"3000";
    tmp(70186) := x"3820";
    tmp(70187) := x"3820";
    tmp(70188) := x"3000";
    tmp(70189) := x"4020";
    tmp(70190) := x"3820";
    tmp(70191) := x"3800";
    tmp(70192) := x"3800";
    tmp(70193) := x"4820";
    tmp(70194) := x"3000";
    tmp(70195) := x"3000";
    tmp(70196) := x"3020";
    tmp(70197) := x"3820";
    tmp(70198) := x"3820";
    tmp(70199) := x"2800";
    tmp(70200) := x"1000";
    tmp(70201) := x"1800";
    tmp(70202) := x"2000";
    tmp(70203) := x"2000";
    tmp(70204) := x"3000";
    tmp(70205) := x"3800";
    tmp(70206) := x"3800";
    tmp(70207) := x"3800";
    tmp(70208) := x"3800";
    tmp(70209) := x"2800";
    tmp(70210) := x"3820";
    tmp(70211) := x"2000";
    tmp(70212) := x"1800";
    tmp(70213) := x"3820";
    tmp(70214) := x"1000";
    tmp(70215) := x"1000";
    tmp(70216) := x"1800";
    tmp(70217) := x"4020";
    tmp(70218) := x"3820";
    tmp(70219) := x"3000";
    tmp(70220) := x"2820";
    tmp(70221) := x"2020";
    tmp(70222) := x"1000";
    tmp(70223) := x"3020";
    tmp(70224) := x"5021";
    tmp(70225) := x"3861";
    tmp(70226) := x"28a1";
    tmp(70227) := x"20a1";
    tmp(70228) := x"18a1";
    tmp(70229) := x"18a1";
    tmp(70230) := x"18a1";
    tmp(70231) := x"18a1";
    tmp(70232) := x"18a1";
    tmp(70233) := x"18a1";
    tmp(70234) := x"1881";
    tmp(70235) := x"1081";
    tmp(70236) := x"1081";
    tmp(70237) := x"1081";
    tmp(70238) := x"1081";
    tmp(70239) := x"1081";
    tmp(70240) := x"1081";
    tmp(70241) := x"1081";
    tmp(70242) := x"1081";
    tmp(70243) := x"1081";
    tmp(70244) := x"1061";
    tmp(70245) := x"1061";
    tmp(70246) := x"1061";
    tmp(70247) := x"1061";
    tmp(70248) := x"1061";
    tmp(70249) := x"0861";
    tmp(70250) := x"0840";
    tmp(70251) := x"0840";
    tmp(70252) := x"0840";
    tmp(70253) := x"0840";
    tmp(70254) := x"0840";
    tmp(70255) := x"0840";
    tmp(70256) := x"0820";
    tmp(70257) := x"0820";
    tmp(70258) := x"0820";
    tmp(70259) := x"0820";
    tmp(70260) := x"0820";
    tmp(70261) := x"0820";
    tmp(70262) := x"0820";
    tmp(70263) := x"0820";
    tmp(70264) := x"0820";
    tmp(70265) := x"0820";
    tmp(70266) := x"0820";
    tmp(70267) := x"0820";
    tmp(70268) := x"0820";
    tmp(70269) := x"0820";
    tmp(70270) := x"0840";
    tmp(70271) := x"0820";
    tmp(70272) := x"0840";
    tmp(70273) := x"0840";
    tmp(70274) := x"0840";
    tmp(70275) := x"0841";
    tmp(70276) := x"0861";
    tmp(70277) := x"1061";
    tmp(70278) := x"1061";
    tmp(70279) := x"1081";
    tmp(70280) := x"10a2";
    tmp(70281) := x"10a2";
    tmp(70282) := x"18a2";
    tmp(70283) := x"18c2";
    tmp(70284) := x"18c2";
    tmp(70285) := x"18e3";
    tmp(70286) := x"2103";
    tmp(70287) := x"2124";
    tmp(70288) := x"2945";
    tmp(70289) := x"3165";
    tmp(70290) := x"31a6";
    tmp(70291) := x"39c7";
    tmp(70292) := x"39e8";
    tmp(70293) := x"4229";
    tmp(70294) := x"4a4a";
    tmp(70295) := x"4a6b";
    tmp(70296) := x"526b";
    tmp(70297) := x"526b";
    tmp(70298) := x"526b";
    tmp(70299) := x"528c";
    tmp(70300) := x"528c";
    tmp(70301) := x"526c";
    tmp(70302) := x"526c";
    tmp(70303) := x"528c";
    tmp(70304) := x"528c";
    tmp(70305) := x"526b";
    tmp(70306) := x"528c";
    tmp(70307) := x"524c";
    tmp(70308) := x"526c";
    tmp(70309) := x"4a6b";
    tmp(70310) := x"4a4b";
    tmp(70311) := x"4a4b";
    tmp(70312) := x"422a";
    tmp(70313) := x"4209";
    tmp(70314) := x"3a09";
    tmp(70315) := x"39c8";
    tmp(70316) := x"31a7";
    tmp(70317) := x"3187";
    tmp(70318) := x"3186";
    tmp(70319) := x"2986";
    tmp(70320) := x"0000";
    tmp(70321) := x"0041";
    tmp(70322) := x"0041";
    tmp(70323) := x"0041";
    tmp(70324) := x"0041";
    tmp(70325) := x"0041";
    tmp(70326) := x"0041";
    tmp(70327) := x"0041";
    tmp(70328) := x"0041";
    tmp(70329) := x"0041";
    tmp(70330) := x"0041";
    tmp(70331) := x"0061";
    tmp(70332) := x"0041";
    tmp(70333) := x"0041";
    tmp(70334) := x"0061";
    tmp(70335) := x"0061";
    tmp(70336) := x"0061";
    tmp(70337) := x"0061";
    tmp(70338) := x"0061";
    tmp(70339) := x"0061";
    tmp(70340) := x"0041";
    tmp(70341) := x"0041";
    tmp(70342) := x"0061";
    tmp(70343) := x"0061";
    tmp(70344) := x"0061";
    tmp(70345) := x"0041";
    tmp(70346) := x"0041";
    tmp(70347) := x"0041";
    tmp(70348) := x"0041";
    tmp(70349) := x"0061";
    tmp(70350) := x"0061";
    tmp(70351) := x"0061";
    tmp(70352) := x"0061";
    tmp(70353) := x"0062";
    tmp(70354) := x"0061";
    tmp(70355) := x"0061";
    tmp(70356) := x"0041";
    tmp(70357) := x"0041";
    tmp(70358) := x"0062";
    tmp(70359) := x"0062";
    tmp(70360) := x"0062";
    tmp(70361) := x"0061";
    tmp(70362) := x"0061";
    tmp(70363) := x"0041";
    tmp(70364) := x"0041";
    tmp(70365) := x"0041";
    tmp(70366) := x"0061";
    tmp(70367) := x"0041";
    tmp(70368) := x"0041";
    tmp(70369) := x"0061";
    tmp(70370) := x"0061";
    tmp(70371) := x"0061";
    tmp(70372) := x"0061";
    tmp(70373) := x"0061";
    tmp(70374) := x"0061";
    tmp(70375) := x"0081";
    tmp(70376) := x"0081";
    tmp(70377) := x"0081";
    tmp(70378) := x"0081";
    tmp(70379) := x"0881";
    tmp(70380) := x"0081";
    tmp(70381) := x"0081";
    tmp(70382) := x"0881";
    tmp(70383) := x"0881";
    tmp(70384) := x"0881";
    tmp(70385) := x"0881";
    tmp(70386) := x"0881";
    tmp(70387) := x"0881";
    tmp(70388) := x"0881";
    tmp(70389) := x"0861";
    tmp(70390) := x"0840";
    tmp(70391) := x"0820";
    tmp(70392) := x"0820";
    tmp(70393) := x"0820";
    tmp(70394) := x"0820";
    tmp(70395) := x"0800";
    tmp(70396) := x"0820";
    tmp(70397) := x"0800";
    tmp(70398) := x"0800";
    tmp(70399) := x"1000";
    tmp(70400) := x"1800";
    tmp(70401) := x"2000";
    tmp(70402) := x"2800";
    tmp(70403) := x"2000";
    tmp(70404) := x"2000";
    tmp(70405) := x"1800";
    tmp(70406) := x"1000";
    tmp(70407) := x"1000";
    tmp(70408) := x"1800";
    tmp(70409) := x"1800";
    tmp(70410) := x"2000";
    tmp(70411) := x"2000";
    tmp(70412) := x"2000";
    tmp(70413) := x"2000";
    tmp(70414) := x"2020";
    tmp(70415) := x"1800";
    tmp(70416) := x"2000";
    tmp(70417) := x"2800";
    tmp(70418) := x"3000";
    tmp(70419) := x"3800";
    tmp(70420) := x"4020";
    tmp(70421) := x"3000";
    tmp(70422) := x"2800";
    tmp(70423) := x"2800";
    tmp(70424) := x"3000";
    tmp(70425) := x"3820";
    tmp(70426) := x"4020";
    tmp(70427) := x"4020";
    tmp(70428) := x"3000";
    tmp(70429) := x"3800";
    tmp(70430) := x"4000";
    tmp(70431) := x"4000";
    tmp(70432) := x"4000";
    tmp(70433) := x"5020";
    tmp(70434) := x"3800";
    tmp(70435) := x"4020";
    tmp(70436) := x"5020";
    tmp(70437) := x"4820";
    tmp(70438) := x"4820";
    tmp(70439) := x"3820";
    tmp(70440) := x"1000";
    tmp(70441) := x"1000";
    tmp(70442) := x"1800";
    tmp(70443) := x"3000";
    tmp(70444) := x"3000";
    tmp(70445) := x"3800";
    tmp(70446) := x"3800";
    tmp(70447) := x"3800";
    tmp(70448) := x"2800";
    tmp(70449) := x"3020";
    tmp(70450) := x"2000";
    tmp(70451) := x"1800";
    tmp(70452) := x"3020";
    tmp(70453) := x"1820";
    tmp(70454) := x"0800";
    tmp(70455) := x"1800";
    tmp(70456) := x"3820";
    tmp(70457) := x"3820";
    tmp(70458) := x"3000";
    tmp(70459) := x"2820";
    tmp(70460) := x"2840";
    tmp(70461) := x"1020";
    tmp(70462) := x"2020";
    tmp(70463) := x"4841";
    tmp(70464) := x"3841";
    tmp(70465) := x"28a1";
    tmp(70466) := x"20a2";
    tmp(70467) := x"18a1";
    tmp(70468) := x"18a1";
    tmp(70469) := x"18a1";
    tmp(70470) := x"18a1";
    tmp(70471) := x"18a1";
    tmp(70472) := x"18a1";
    tmp(70473) := x"18a1";
    tmp(70474) := x"1081";
    tmp(70475) := x"1081";
    tmp(70476) := x"1081";
    tmp(70477) := x"1081";
    tmp(70478) := x"1081";
    tmp(70479) := x"1081";
    tmp(70480) := x"1081";
    tmp(70481) := x"1061";
    tmp(70482) := x"1061";
    tmp(70483) := x"1061";
    tmp(70484) := x"1061";
    tmp(70485) := x"1061";
    tmp(70486) := x"0861";
    tmp(70487) := x"1061";
    tmp(70488) := x"0860";
    tmp(70489) := x"0840";
    tmp(70490) := x"0840";
    tmp(70491) := x"0840";
    tmp(70492) := x"0840";
    tmp(70493) := x"0840";
    tmp(70494) := x"0840";
    tmp(70495) := x"0820";
    tmp(70496) := x"0820";
    tmp(70497) := x"0820";
    tmp(70498) := x"0820";
    tmp(70499) := x"0820";
    tmp(70500) := x"0820";
    tmp(70501) := x"0820";
    tmp(70502) := x"0820";
    tmp(70503) := x"0820";
    tmp(70504) := x"0820";
    tmp(70505) := x"0820";
    tmp(70506) := x"0820";
    tmp(70507) := x"0820";
    tmp(70508) := x"0820";
    tmp(70509) := x"0820";
    tmp(70510) := x"0820";
    tmp(70511) := x"0820";
    tmp(70512) := x"0820";
    tmp(70513) := x"0820";
    tmp(70514) := x"0820";
    tmp(70515) := x"0840";
    tmp(70516) := x"0840";
    tmp(70517) := x"0841";
    tmp(70518) := x"0861";
    tmp(70519) := x"1061";
    tmp(70520) := x"1081";
    tmp(70521) := x"1081";
    tmp(70522) := x"10a2";
    tmp(70523) := x"10a2";
    tmp(70524) := x"10c2";
    tmp(70525) := x"18c2";
    tmp(70526) := x"18e3";
    tmp(70527) := x"2103";
    tmp(70528) := x"2104";
    tmp(70529) := x"2924";
    tmp(70530) := x"2965";
    tmp(70531) := x"3165";
    tmp(70532) := x"31a6";
    tmp(70533) := x"39c7";
    tmp(70534) := x"41e8";
    tmp(70535) := x"4209";
    tmp(70536) := x"422a";
    tmp(70537) := x"4a2a";
    tmp(70538) := x"422a";
    tmp(70539) := x"4a2a";
    tmp(70540) := x"4a2a";
    tmp(70541) := x"4a4b";
    tmp(70542) := x"4a4b";
    tmp(70543) := x"4a4b";
    tmp(70544) := x"4a4b";
    tmp(70545) := x"4a4a";
    tmp(70546) := x"4a4a";
    tmp(70547) := x"4a2a";
    tmp(70548) := x"422a";
    tmp(70549) := x"422a";
    tmp(70550) := x"422a";
    tmp(70551) := x"4209";
    tmp(70552) := x"39e8";
    tmp(70553) := x"39c8";
    tmp(70554) := x"39c7";
    tmp(70555) := x"31a7";
    tmp(70556) := x"2986";
    tmp(70557) := x"2966";
    tmp(70558) := x"2965";
    tmp(70559) := x"2945";
    tmp(70560) := x"0000";
    tmp(70561) := x"0020";
    tmp(70562) := x"0021";
    tmp(70563) := x"0041";
    tmp(70564) := x"0041";
    tmp(70565) := x"0041";
    tmp(70566) := x"0041";
    tmp(70567) := x"0041";
    tmp(70568) := x"0041";
    tmp(70569) := x"0041";
    tmp(70570) := x"0061";
    tmp(70571) := x"0041";
    tmp(70572) := x"0061";
    tmp(70573) := x"0061";
    tmp(70574) := x"0061";
    tmp(70575) := x"0061";
    tmp(70576) := x"0061";
    tmp(70577) := x"0061";
    tmp(70578) := x"0062";
    tmp(70579) := x"0062";
    tmp(70580) := x"0062";
    tmp(70581) := x"0062";
    tmp(70582) := x"0061";
    tmp(70583) := x"0061";
    tmp(70584) := x"0061";
    tmp(70585) := x"0041";
    tmp(70586) := x"0041";
    tmp(70587) := x"0041";
    tmp(70588) := x"0041";
    tmp(70589) := x"0041";
    tmp(70590) := x"0041";
    tmp(70591) := x"0041";
    tmp(70592) := x"0061";
    tmp(70593) := x"0061";
    tmp(70594) := x"0061";
    tmp(70595) := x"0061";
    tmp(70596) := x"0061";
    tmp(70597) := x"0061";
    tmp(70598) := x"0061";
    tmp(70599) := x"0061";
    tmp(70600) := x"0061";
    tmp(70601) := x"0061";
    tmp(70602) := x"0061";
    tmp(70603) := x"0041";
    tmp(70604) := x"0041";
    tmp(70605) := x"0021";
    tmp(70606) := x"0041";
    tmp(70607) := x"0041";
    tmp(70608) := x"0041";
    tmp(70609) := x"0061";
    tmp(70610) := x"0061";
    tmp(70611) := x"0061";
    tmp(70612) := x"0061";
    tmp(70613) := x"0061";
    tmp(70614) := x"0061";
    tmp(70615) := x"0061";
    tmp(70616) := x"0061";
    tmp(70617) := x"0061";
    tmp(70618) := x"0061";
    tmp(70619) := x"0061";
    tmp(70620) := x"0061";
    tmp(70621) := x"0060";
    tmp(70622) := x"0060";
    tmp(70623) := x"0060";
    tmp(70624) := x"0060";
    tmp(70625) := x"0040";
    tmp(70626) := x"0040";
    tmp(70627) := x"0040";
    tmp(70628) := x"0040";
    tmp(70629) := x"0040";
    tmp(70630) := x"0020";
    tmp(70631) := x"0820";
    tmp(70632) := x"0820";
    tmp(70633) := x"0820";
    tmp(70634) := x"0800";
    tmp(70635) := x"0820";
    tmp(70636) := x"0820";
    tmp(70637) := x"0820";
    tmp(70638) := x"0820";
    tmp(70639) := x"0800";
    tmp(70640) := x"1000";
    tmp(70641) := x"1800";
    tmp(70642) := x"2000";
    tmp(70643) := x"2800";
    tmp(70644) := x"2000";
    tmp(70645) := x"1000";
    tmp(70646) := x"1000";
    tmp(70647) := x"1000";
    tmp(70648) := x"1000";
    tmp(70649) := x"1800";
    tmp(70650) := x"1800";
    tmp(70651) := x"1800";
    tmp(70652) := x"2000";
    tmp(70653) := x"2000";
    tmp(70654) := x"2000";
    tmp(70655) := x"1800";
    tmp(70656) := x"2000";
    tmp(70657) := x"2000";
    tmp(70658) := x"2800";
    tmp(70659) := x"3000";
    tmp(70660) := x"3800";
    tmp(70661) := x"3000";
    tmp(70662) := x"2800";
    tmp(70663) := x"2800";
    tmp(70664) := x"3820";
    tmp(70665) := x"3820";
    tmp(70666) := x"3820";
    tmp(70667) := x"3820";
    tmp(70668) := x"3800";
    tmp(70669) := x"4000";
    tmp(70670) := x"4800";
    tmp(70671) := x"5000";
    tmp(70672) := x"4800";
    tmp(70673) := x"5020";
    tmp(70674) := x"4020";
    tmp(70675) := x"3000";
    tmp(70676) := x"4020";
    tmp(70677) := x"5020";
    tmp(70678) := x"4020";
    tmp(70679) := x"4020";
    tmp(70680) := x"1800";
    tmp(70681) := x"2000";
    tmp(70682) := x"2800";
    tmp(70683) := x"3000";
    tmp(70684) := x"3000";
    tmp(70685) := x"3800";
    tmp(70686) := x"3800";
    tmp(70687) := x"3000";
    tmp(70688) := x"3820";
    tmp(70689) := x"2800";
    tmp(70690) := x"2000";
    tmp(70691) := x"4020";
    tmp(70692) := x"2020";
    tmp(70693) := x"1840";
    tmp(70694) := x"1820";
    tmp(70695) := x"3020";
    tmp(70696) := x"4020";
    tmp(70697) := x"3000";
    tmp(70698) := x"2800";
    tmp(70699) := x"2861";
    tmp(70700) := x"1840";
    tmp(70701) := x"1820";
    tmp(70702) := x"3841";
    tmp(70703) := x"3841";
    tmp(70704) := x"2881";
    tmp(70705) := x"20a2";
    tmp(70706) := x"18a2";
    tmp(70707) := x"18a1";
    tmp(70708) := x"18a1";
    tmp(70709) := x"18a1";
    tmp(70710) := x"18a1";
    tmp(70711) := x"18a1";
    tmp(70712) := x"10a1";
    tmp(70713) := x"1081";
    tmp(70714) := x"1081";
    tmp(70715) := x"1081";
    tmp(70716) := x"1081";
    tmp(70717) := x"1081";
    tmp(70718) := x"1081";
    tmp(70719) := x"1061";
    tmp(70720) := x"1061";
    tmp(70721) := x"1061";
    tmp(70722) := x"1061";
    tmp(70723) := x"1061";
    tmp(70724) := x"1061";
    tmp(70725) := x"0860";
    tmp(70726) := x"0860";
    tmp(70727) := x"0840";
    tmp(70728) := x"0840";
    tmp(70729) := x"0840";
    tmp(70730) := x"0840";
    tmp(70731) := x"0840";
    tmp(70732) := x"0840";
    tmp(70733) := x"0820";
    tmp(70734) := x"0820";
    tmp(70735) := x"0820";
    tmp(70736) := x"0820";
    tmp(70737) := x"0820";
    tmp(70738) := x"0820";
    tmp(70739) := x"0820";
    tmp(70740) := x"0820";
    tmp(70741) := x"0820";
    tmp(70742) := x"0820";
    tmp(70743) := x"0820";
    tmp(70744) := x"0820";
    tmp(70745) := x"0820";
    tmp(70746) := x"0820";
    tmp(70747) := x"0820";
    tmp(70748) := x"0820";
    tmp(70749) := x"0820";
    tmp(70750) := x"0820";
    tmp(70751) := x"0820";
    tmp(70752) := x"0820";
    tmp(70753) := x"0820";
    tmp(70754) := x"0820";
    tmp(70755) := x"0820";
    tmp(70756) := x"0840";
    tmp(70757) := x"0840";
    tmp(70758) := x"0841";
    tmp(70759) := x"0861";
    tmp(70760) := x"0861";
    tmp(70761) := x"1061";
    tmp(70762) := x"1081";
    tmp(70763) := x"1081";
    tmp(70764) := x"10a2";
    tmp(70765) := x"10a2";
    tmp(70766) := x"18c2";
    tmp(70767) := x"18c3";
    tmp(70768) := x"1903";
    tmp(70769) := x"2104";
    tmp(70770) := x"2124";
    tmp(70771) := x"2965";
    tmp(70772) := x"2965";
    tmp(70773) := x"3185";
    tmp(70774) := x"31a6";
    tmp(70775) := x"39a7";
    tmp(70776) := x"39c7";
    tmp(70777) := x"39e8";
    tmp(70778) := x"41e9";
    tmp(70779) := x"41e8";
    tmp(70780) := x"4209";
    tmp(70781) := x"4209";
    tmp(70782) := x"4209";
    tmp(70783) := x"420a";
    tmp(70784) := x"4209";
    tmp(70785) := x"4209";
    tmp(70786) := x"4209";
    tmp(70787) := x"39e9";
    tmp(70788) := x"39e8";
    tmp(70789) := x"4208";
    tmp(70790) := x"39c7";
    tmp(70791) := x"31a7";
    tmp(70792) := x"31a7";
    tmp(70793) := x"3186";
    tmp(70794) := x"2986";
    tmp(70795) := x"2966";
    tmp(70796) := x"2965";
    tmp(70797) := x"2145";
    tmp(70798) := x"2144";
    tmp(70799) := x"2104";
    tmp(70800) := x"0000";
    tmp(70801) := x"0000";
    tmp(70802) := x"0000";
    tmp(70803) := x"0020";
    tmp(70804) := x"0020";
    tmp(70805) := x"0021";
    tmp(70806) := x"0041";
    tmp(70807) := x"0041";
    tmp(70808) := x"0041";
    tmp(70809) := x"0041";
    tmp(70810) := x"0041";
    tmp(70811) := x"0061";
    tmp(70812) := x"0061";
    tmp(70813) := x"0061";
    tmp(70814) := x"0061";
    tmp(70815) := x"0061";
    tmp(70816) := x"0062";
    tmp(70817) := x"0061";
    tmp(70818) := x"0061";
    tmp(70819) := x"0062";
    tmp(70820) := x"0062";
    tmp(70821) := x"0062";
    tmp(70822) := x"0062";
    tmp(70823) := x"0061";
    tmp(70824) := x"0041";
    tmp(70825) := x"0020";
    tmp(70826) := x"0021";
    tmp(70827) := x"0041";
    tmp(70828) := x"0041";
    tmp(70829) := x"0041";
    tmp(70830) := x"0041";
    tmp(70831) := x"0041";
    tmp(70832) := x"0041";
    tmp(70833) := x"0041";
    tmp(70834) := x"0061";
    tmp(70835) := x"0061";
    tmp(70836) := x"0041";
    tmp(70837) := x"0041";
    tmp(70838) := x"0061";
    tmp(70839) := x"0061";
    tmp(70840) := x"0061";
    tmp(70841) := x"0041";
    tmp(70842) := x"0041";
    tmp(70843) := x"0041";
    tmp(70844) := x"0041";
    tmp(70845) := x"0061";
    tmp(70846) := x"0041";
    tmp(70847) := x"0040";
    tmp(70848) := x"0040";
    tmp(70849) := x"0061";
    tmp(70850) := x"0061";
    tmp(70851) := x"0061";
    tmp(70852) := x"0061";
    tmp(70853) := x"0061";
    tmp(70854) := x"0061";
    tmp(70855) := x"0060";
    tmp(70856) := x"0060";
    tmp(70857) := x"0060";
    tmp(70858) := x"0060";
    tmp(70859) := x"0860";
    tmp(70860) := x"0860";
    tmp(70861) := x"0860";
    tmp(70862) := x"0880";
    tmp(70863) := x"0880";
    tmp(70864) := x"0880";
    tmp(70865) := x"0880";
    tmp(70866) := x"0880";
    tmp(70867) := x"0881";
    tmp(70868) := x"0881";
    tmp(70869) := x"0881";
    tmp(70870) := x"0881";
    tmp(70871) := x"0861";
    tmp(70872) := x"0861";
    tmp(70873) := x"0841";
    tmp(70874) := x"0820";
    tmp(70875) := x"0820";
    tmp(70876) := x"0820";
    tmp(70877) := x"0820";
    tmp(70878) := x"0820";
    tmp(70879) := x"0820";
    tmp(70880) := x"0800";
    tmp(70881) := x"1000";
    tmp(70882) := x"1800";
    tmp(70883) := x"2000";
    tmp(70884) := x"1000";
    tmp(70885) := x"0800";
    tmp(70886) := x"1000";
    tmp(70887) := x"1000";
    tmp(70888) := x"1000";
    tmp(70889) := x"1800";
    tmp(70890) := x"1800";
    tmp(70891) := x"1800";
    tmp(70892) := x"2000";
    tmp(70893) := x"2000";
    tmp(70894) := x"2020";
    tmp(70895) := x"2020";
    tmp(70896) := x"2000";
    tmp(70897) := x"2000";
    tmp(70898) := x"2800";
    tmp(70899) := x"3000";
    tmp(70900) := x"3000";
    tmp(70901) := x"2800";
    tmp(70902) := x"2800";
    tmp(70903) := x"3000";
    tmp(70904) := x"3020";
    tmp(70905) := x"3820";
    tmp(70906) := x"4020";
    tmp(70907) := x"5020";
    tmp(70908) := x"5020";
    tmp(70909) := x"4820";
    tmp(70910) := x"4800";
    tmp(70911) := x"5020";
    tmp(70912) := x"4800";
    tmp(70913) := x"4820";
    tmp(70914) := x"4020";
    tmp(70915) := x"4020";
    tmp(70916) := x"5020";
    tmp(70917) := x"4820";
    tmp(70918) := x"4820";
    tmp(70919) := x"4820";
    tmp(70920) := x"1800";
    tmp(70921) := x"3820";
    tmp(70922) := x"3000";
    tmp(70923) := x"3000";
    tmp(70924) := x"3000";
    tmp(70925) := x"3000";
    tmp(70926) := x"3000";
    tmp(70927) := x"3000";
    tmp(70928) := x"2800";
    tmp(70929) := x"2800";
    tmp(70930) := x"4020";
    tmp(70931) := x"2020";
    tmp(70932) := x"1840";
    tmp(70933) := x"2881";
    tmp(70934) := x"2020";
    tmp(70935) := x"2000";
    tmp(70936) := x"3020";
    tmp(70937) := x"2820";
    tmp(70938) := x"3081";
    tmp(70939) := x"2061";
    tmp(70940) := x"1020";
    tmp(70941) := x"2861";
    tmp(70942) := x"3081";
    tmp(70943) := x"2881";
    tmp(70944) := x"20c2";
    tmp(70945) := x"18c2";
    tmp(70946) := x"18a1";
    tmp(70947) := x"18a1";
    tmp(70948) := x"18a1";
    tmp(70949) := x"10a1";
    tmp(70950) := x"18a1";
    tmp(70951) := x"18a1";
    tmp(70952) := x"1081";
    tmp(70953) := x"1081";
    tmp(70954) := x"1081";
    tmp(70955) := x"1081";
    tmp(70956) := x"1081";
    tmp(70957) := x"1081";
    tmp(70958) := x"1061";
    tmp(70959) := x"1061";
    tmp(70960) := x"1061";
    tmp(70961) := x"1061";
    tmp(70962) := x"0860";
    tmp(70963) := x"0861";
    tmp(70964) := x"0860";
    tmp(70965) := x"0840";
    tmp(70966) := x"0840";
    tmp(70967) := x"0840";
    tmp(70968) := x"0840";
    tmp(70969) := x"0840";
    tmp(70970) := x"0840";
    tmp(70971) := x"0840";
    tmp(70972) := x"0820";
    tmp(70973) := x"0820";
    tmp(70974) := x"0820";
    tmp(70975) := x"0820";
    tmp(70976) := x"0820";
    tmp(70977) := x"0820";
    tmp(70978) := x"0820";
    tmp(70979) := x"0820";
    tmp(70980) := x"0820";
    tmp(70981) := x"0820";
    tmp(70982) := x"0820";
    tmp(70983) := x"0820";
    tmp(70984) := x"0820";
    tmp(70985) := x"0820";
    tmp(70986) := x"0820";
    tmp(70987) := x"0020";
    tmp(70988) := x"0020";
    tmp(70989) := x"0020";
    tmp(70990) := x"0020";
    tmp(70991) := x"0020";
    tmp(70992) := x"0020";
    tmp(70993) := x"0820";
    tmp(70994) := x"0820";
    tmp(70995) := x"0820";
    tmp(70996) := x"0820";
    tmp(70997) := x"0820";
    tmp(70998) := x"0840";
    tmp(70999) := x"0840";
    tmp(71000) := x"0841";
    tmp(71001) := x"0861";
    tmp(71002) := x"0861";
    tmp(71003) := x"0861";
    tmp(71004) := x"1081";
    tmp(71005) := x"1081";
    tmp(71006) := x"10a2";
    tmp(71007) := x"10a2";
    tmp(71008) := x"18c2";
    tmp(71009) := x"18e3";
    tmp(71010) := x"18e3";
    tmp(71011) := x"2104";
    tmp(71012) := x"2124";
    tmp(71013) := x"2945";
    tmp(71014) := x"2965";
    tmp(71015) := x"2965";
    tmp(71016) := x"3186";
    tmp(71017) := x"3186";
    tmp(71018) := x"31a7";
    tmp(71019) := x"39a7";
    tmp(71020) := x"39c7";
    tmp(71021) := x"39c7";
    tmp(71022) := x"39c7";
    tmp(71023) := x"39c7";
    tmp(71024) := x"39c8";
    tmp(71025) := x"39c7";
    tmp(71026) := x"39c7";
    tmp(71027) := x"31c7";
    tmp(71028) := x"31c7";
    tmp(71029) := x"3186";
    tmp(71030) := x"2986";
    tmp(71031) := x"2965";
    tmp(71032) := x"2945";
    tmp(71033) := x"2945";
    tmp(71034) := x"2145";
    tmp(71035) := x"2124";
    tmp(71036) := x"2124";
    tmp(71037) := x"1904";
    tmp(71038) := x"1903";
    tmp(71039) := x"18e3";
    tmp(71040) := x"0000";
    tmp(71041) := x"0021";
    tmp(71042) := x"0020";
    tmp(71043) := x"0020";
    tmp(71044) := x"0000";
    tmp(71045) := x"0000";
    tmp(71046) := x"0020";
    tmp(71047) := x"0020";
    tmp(71048) := x"0021";
    tmp(71049) := x"0021";
    tmp(71050) := x"0041";
    tmp(71051) := x"0041";
    tmp(71052) := x"0041";
    tmp(71053) := x"0041";
    tmp(71054) := x"0061";
    tmp(71055) := x"0061";
    tmp(71056) := x"0062";
    tmp(71057) := x"0061";
    tmp(71058) := x"0061";
    tmp(71059) := x"0062";
    tmp(71060) := x"0062";
    tmp(71061) := x"0062";
    tmp(71062) := x"0061";
    tmp(71063) := x"0041";
    tmp(71064) := x"0020";
    tmp(71065) := x"0020";
    tmp(71066) := x"0021";
    tmp(71067) := x"0041";
    tmp(71068) := x"0041";
    tmp(71069) := x"0041";
    tmp(71070) := x"0041";
    tmp(71071) := x"0041";
    tmp(71072) := x"0041";
    tmp(71073) := x"0041";
    tmp(71074) := x"0061";
    tmp(71075) := x"0061";
    tmp(71076) := x"0061";
    tmp(71077) := x"0061";
    tmp(71078) := x"0061";
    tmp(71079) := x"0061";
    tmp(71080) := x"0061";
    tmp(71081) := x"0041";
    tmp(71082) := x"0041";
    tmp(71083) := x"0040";
    tmp(71084) := x"0040";
    tmp(71085) := x"0041";
    tmp(71086) := x"0040";
    tmp(71087) := x"0020";
    tmp(71088) := x"0020";
    tmp(71089) := x"0040";
    tmp(71090) := x"0040";
    tmp(71091) := x"0040";
    tmp(71092) := x"0040";
    tmp(71093) := x"0040";
    tmp(71094) := x"0040";
    tmp(71095) := x"0040";
    tmp(71096) := x"0060";
    tmp(71097) := x"0060";
    tmp(71098) := x"0060";
    tmp(71099) := x"0040";
    tmp(71100) := x"0060";
    tmp(71101) := x"0060";
    tmp(71102) := x"0060";
    tmp(71103) := x"0060";
    tmp(71104) := x"0060";
    tmp(71105) := x"0060";
    tmp(71106) := x"0040";
    tmp(71107) := x"0040";
    tmp(71108) := x"0860";
    tmp(71109) := x"0860";
    tmp(71110) := x"0061";
    tmp(71111) := x"0061";
    tmp(71112) := x"0061";
    tmp(71113) := x"0061";
    tmp(71114) := x"0861";
    tmp(71115) := x"0861";
    tmp(71116) := x"0841";
    tmp(71117) := x"0841";
    tmp(71118) := x"0820";
    tmp(71119) := x"0820";
    tmp(71120) := x"0820";
    tmp(71121) := x"0820";
    tmp(71122) := x"0800";
    tmp(71123) := x"1000";
    tmp(71124) := x"0800";
    tmp(71125) := x"0800";
    tmp(71126) := x"1000";
    tmp(71127) := x"1000";
    tmp(71128) := x"1800";
    tmp(71129) := x"1800";
    tmp(71130) := x"1800";
    tmp(71131) := x"1800";
    tmp(71132) := x"2000";
    tmp(71133) := x"2000";
    tmp(71134) := x"2000";
    tmp(71135) := x"2820";
    tmp(71136) := x"2020";
    tmp(71137) := x"2000";
    tmp(71138) := x"2000";
    tmp(71139) := x"2800";
    tmp(71140) := x"2800";
    tmp(71141) := x"2800";
    tmp(71142) := x"2800";
    tmp(71143) := x"3020";
    tmp(71144) := x"3020";
    tmp(71145) := x"4840";
    tmp(71146) := x"5861";
    tmp(71147) := x"5840";
    tmp(71148) := x"5040";
    tmp(71149) := x"4820";
    tmp(71150) := x"5020";
    tmp(71151) := x"5820";
    tmp(71152) := x"5020";
    tmp(71153) := x"4020";
    tmp(71154) := x"4020";
    tmp(71155) := x"4820";
    tmp(71156) := x"5020";
    tmp(71157) := x"4020";
    tmp(71158) := x"4020";
    tmp(71159) := x"4020";
    tmp(71160) := x"3820";
    tmp(71161) := x"3820";
    tmp(71162) := x"3000";
    tmp(71163) := x"3000";
    tmp(71164) := x"3800";
    tmp(71165) := x"3800";
    tmp(71166) := x"3000";
    tmp(71167) := x"3000";
    tmp(71168) := x"2800";
    tmp(71169) := x"3820";
    tmp(71170) := x"2820";
    tmp(71171) := x"1820";
    tmp(71172) := x"20c2";
    tmp(71173) := x"2861";
    tmp(71174) := x"2020";
    tmp(71175) := x"3841";
    tmp(71176) := x"3041";
    tmp(71177) := x"2881";
    tmp(71178) := x"20a1";
    tmp(71179) := x"1841";
    tmp(71180) := x"1861";
    tmp(71181) := x"28a2";
    tmp(71182) := x"20a2";
    tmp(71183) := x"20a2";
    tmp(71184) := x"18a2";
    tmp(71185) := x"18a1";
    tmp(71186) := x"18a1";
    tmp(71187) := x"18a1";
    tmp(71188) := x"18a1";
    tmp(71189) := x"18a1";
    tmp(71190) := x"1081";
    tmp(71191) := x"1081";
    tmp(71192) := x"1081";
    tmp(71193) := x"1081";
    tmp(71194) := x"1081";
    tmp(71195) := x"1081";
    tmp(71196) := x"1061";
    tmp(71197) := x"1061";
    tmp(71198) := x"1061";
    tmp(71199) := x"1061";
    tmp(71200) := x"1061";
    tmp(71201) := x"0861";
    tmp(71202) := x"0840";
    tmp(71203) := x"0840";
    tmp(71204) := x"0840";
    tmp(71205) := x"0840";
    tmp(71206) := x"0840";
    tmp(71207) := x"0840";
    tmp(71208) := x"0840";
    tmp(71209) := x"0840";
    tmp(71210) := x"0820";
    tmp(71211) := x"0820";
    tmp(71212) := x"0820";
    tmp(71213) := x"0820";
    tmp(71214) := x"0820";
    tmp(71215) := x"0820";
    tmp(71216) := x"0820";
    tmp(71217) := x"0820";
    tmp(71218) := x"0820";
    tmp(71219) := x"0820";
    tmp(71220) := x"0820";
    tmp(71221) := x"0820";
    tmp(71222) := x"0820";
    tmp(71223) := x"0820";
    tmp(71224) := x"0820";
    tmp(71225) := x"0020";
    tmp(71226) := x"0020";
    tmp(71227) := x"0020";
    tmp(71228) := x"0020";
    tmp(71229) := x"0020";
    tmp(71230) := x"0020";
    tmp(71231) := x"0020";
    tmp(71232) := x"0020";
    tmp(71233) := x"0020";
    tmp(71234) := x"0020";
    tmp(71235) := x"0820";
    tmp(71236) := x"0820";
    tmp(71237) := x"0820";
    tmp(71238) := x"0820";
    tmp(71239) := x"0820";
    tmp(71240) := x"0840";
    tmp(71241) := x"0840";
    tmp(71242) := x"0841";
    tmp(71243) := x"0841";
    tmp(71244) := x"0861";
    tmp(71245) := x"1061";
    tmp(71246) := x"1081";
    tmp(71247) := x"1081";
    tmp(71248) := x"10a2";
    tmp(71249) := x"10a2";
    tmp(71250) := x"18c2";
    tmp(71251) := x"18e3";
    tmp(71252) := x"2103";
    tmp(71253) := x"2104";
    tmp(71254) := x"2124";
    tmp(71255) := x"2924";
    tmp(71256) := x"2925";
    tmp(71257) := x"2945";
    tmp(71258) := x"2965";
    tmp(71259) := x"2965";
    tmp(71260) := x"2966";
    tmp(71261) := x"3186";
    tmp(71262) := x"3186";
    tmp(71263) := x"3186";
    tmp(71264) := x"3186";
    tmp(71265) := x"2986";
    tmp(71266) := x"2965";
    tmp(71267) := x"2965";
    tmp(71268) := x"2945";
    tmp(71269) := x"2945";
    tmp(71270) := x"2145";
    tmp(71271) := x"2124";
    tmp(71272) := x"2124";
    tmp(71273) := x"2104";
    tmp(71274) := x"2104";
    tmp(71275) := x"1903";
    tmp(71276) := x"18e3";
    tmp(71277) := x"18e3";
    tmp(71278) := x"18c2";
    tmp(71279) := x"10c2";
    tmp(71280) := x"0000";
    tmp(71281) := x"0021";
    tmp(71282) := x"0021";
    tmp(71283) := x"0021";
    tmp(71284) := x"0041";
    tmp(71285) := x"0041";
    tmp(71286) := x"0021";
    tmp(71287) := x"0021";
    tmp(71288) := x"0021";
    tmp(71289) := x"0021";
    tmp(71290) := x"0021";
    tmp(71291) := x"0021";
    tmp(71292) := x"0041";
    tmp(71293) := x"0041";
    tmp(71294) := x"0041";
    tmp(71295) := x"0041";
    tmp(71296) := x"0041";
    tmp(71297) := x"0061";
    tmp(71298) := x"0061";
    tmp(71299) := x"0061";
    tmp(71300) := x"0062";
    tmp(71301) := x"0061";
    tmp(71302) := x"0041";
    tmp(71303) := x"0021";
    tmp(71304) := x"0020";
    tmp(71305) := x"0020";
    tmp(71306) := x"0021";
    tmp(71307) := x"0041";
    tmp(71308) := x"0041";
    tmp(71309) := x"0041";
    tmp(71310) := x"0041";
    tmp(71311) := x"0041";
    tmp(71312) := x"0041";
    tmp(71313) := x"0041";
    tmp(71314) := x"0061";
    tmp(71315) := x"0061";
    tmp(71316) := x"0061";
    tmp(71317) := x"0061";
    tmp(71318) := x"0061";
    tmp(71319) := x"0061";
    tmp(71320) := x"0061";
    tmp(71321) := x"0041";
    tmp(71322) := x"0040";
    tmp(71323) := x"0040";
    tmp(71324) := x"0040";
    tmp(71325) := x"0040";
    tmp(71326) := x"0040";
    tmp(71327) := x"0020";
    tmp(71328) := x"0020";
    tmp(71329) := x"0040";
    tmp(71330) := x"0040";
    tmp(71331) := x"0040";
    tmp(71332) := x"0040";
    tmp(71333) := x"0040";
    tmp(71334) := x"0040";
    tmp(71335) := x"0040";
    tmp(71336) := x"0040";
    tmp(71337) := x"0040";
    tmp(71338) := x"0040";
    tmp(71339) := x"0040";
    tmp(71340) := x"0040";
    tmp(71341) := x"0040";
    tmp(71342) := x"0040";
    tmp(71343) := x"0040";
    tmp(71344) := x"0040";
    tmp(71345) := x"0040";
    tmp(71346) := x"0040";
    tmp(71347) := x"0040";
    tmp(71348) := x"0060";
    tmp(71349) := x"0060";
    tmp(71350) := x"0061";
    tmp(71351) := x"0061";
    tmp(71352) := x"0061";
    tmp(71353) := x"0061";
    tmp(71354) := x"0061";
    tmp(71355) := x"0861";
    tmp(71356) := x"0861";
    tmp(71357) := x"0840";
    tmp(71358) := x"0840";
    tmp(71359) := x"0820";
    tmp(71360) := x"0840";
    tmp(71361) := x"0840";
    tmp(71362) := x"0820";
    tmp(71363) := x"0820";
    tmp(71364) := x"0800";
    tmp(71365) := x"0800";
    tmp(71366) := x"1000";
    tmp(71367) := x"1800";
    tmp(71368) := x"1800";
    tmp(71369) := x"1800";
    tmp(71370) := x"1800";
    tmp(71371) := x"1800";
    tmp(71372) := x"2000";
    tmp(71373) := x"2000";
    tmp(71374) := x"2000";
    tmp(71375) := x"2820";
    tmp(71376) := x"2020";
    tmp(71377) := x"2020";
    tmp(71378) := x"1800";
    tmp(71379) := x"2000";
    tmp(71380) := x"3020";
    tmp(71381) := x"3820";
    tmp(71382) := x"4820";
    tmp(71383) := x"5040";
    tmp(71384) := x"5040";
    tmp(71385) := x"5040";
    tmp(71386) := x"4840";
    tmp(71387) := x"3820";
    tmp(71388) := x"3820";
    tmp(71389) := x"4020";
    tmp(71390) := x"5020";
    tmp(71391) := x"5020";
    tmp(71392) := x"4820";
    tmp(71393) := x"4000";
    tmp(71394) := x"4820";
    tmp(71395) := x"4020";
    tmp(71396) := x"3800";
    tmp(71397) := x"3800";
    tmp(71398) := x"4020";
    tmp(71399) := x"4820";
    tmp(71400) := x"5840";
    tmp(71401) := x"3000";
    tmp(71402) := x"2800";
    tmp(71403) := x"3000";
    tmp(71404) := x"3800";
    tmp(71405) := x"3000";
    tmp(71406) := x"3000";
    tmp(71407) := x"3000";
    tmp(71408) := x"3000";
    tmp(71409) := x"3020";
    tmp(71410) := x"1820";
    tmp(71411) := x"2081";
    tmp(71412) := x"20c2";
    tmp(71413) := x"2061";
    tmp(71414) := x"2861";
    tmp(71415) := x"2881";
    tmp(71416) := x"28a2";
    tmp(71417) := x"18c2";
    tmp(71418) := x"20a2";
    tmp(71419) := x"20a1";
    tmp(71420) := x"20c2";
    tmp(71421) := x"18c2";
    tmp(71422) := x"18c2";
    tmp(71423) := x"18c2";
    tmp(71424) := x"18a1";
    tmp(71425) := x"18a1";
    tmp(71426) := x"18a1";
    tmp(71427) := x"18a1";
    tmp(71428) := x"10a1";
    tmp(71429) := x"18a1";
    tmp(71430) := x"1081";
    tmp(71431) := x"1081";
    tmp(71432) := x"1081";
    tmp(71433) := x"1081";
    tmp(71434) := x"1081";
    tmp(71435) := x"1061";
    tmp(71436) := x"1061";
    tmp(71437) := x"1061";
    tmp(71438) := x"1061";
    tmp(71439) := x"1061";
    tmp(71440) := x"0861";
    tmp(71441) := x"0840";
    tmp(71442) := x"0840";
    tmp(71443) := x"0840";
    tmp(71444) := x"0840";
    tmp(71445) := x"0840";
    tmp(71446) := x"0840";
    tmp(71447) := x"0840";
    tmp(71448) := x"0840";
    tmp(71449) := x"0820";
    tmp(71450) := x"0820";
    tmp(71451) := x"0820";
    tmp(71452) := x"0820";
    tmp(71453) := x"0820";
    tmp(71454) := x"0820";
    tmp(71455) := x"0820";
    tmp(71456) := x"0820";
    tmp(71457) := x"0820";
    tmp(71458) := x"0820";
    tmp(71459) := x"0820";
    tmp(71460) := x"0020";
    tmp(71461) := x"0020";
    tmp(71462) := x"0020";
    tmp(71463) := x"0020";
    tmp(71464) := x"0020";
    tmp(71465) := x"0020";
    tmp(71466) := x"0020";
    tmp(71467) := x"0020";
    tmp(71468) := x"0020";
    tmp(71469) := x"0020";
    tmp(71470) := x"0020";
    tmp(71471) := x"0020";
    tmp(71472) := x"0020";
    tmp(71473) := x"0020";
    tmp(71474) := x"0020";
    tmp(71475) := x"0020";
    tmp(71476) := x"0020";
    tmp(71477) := x"0820";
    tmp(71478) := x"0820";
    tmp(71479) := x"0820";
    tmp(71480) := x"0820";
    tmp(71481) := x"0820";
    tmp(71482) := x"0840";
    tmp(71483) := x"0840";
    tmp(71484) := x"0841";
    tmp(71485) := x"0841";
    tmp(71486) := x"0861";
    tmp(71487) := x"0861";
    tmp(71488) := x"1081";
    tmp(71489) := x"10a1";
    tmp(71490) := x"10a2";
    tmp(71491) := x"10a2";
    tmp(71492) := x"18c2";
    tmp(71493) := x"18e3";
    tmp(71494) := x"18e3";
    tmp(71495) := x"20e3";
    tmp(71496) := x"2104";
    tmp(71497) := x"2104";
    tmp(71498) := x"2124";
    tmp(71499) := x"2124";
    tmp(71500) := x"2124";
    tmp(71501) := x"2124";
    tmp(71502) := x"2144";
    tmp(71503) := x"2924";
    tmp(71504) := x"2124";
    tmp(71505) := x"2124";
    tmp(71506) := x"2124";
    tmp(71507) := x"2104";
    tmp(71508) := x"2104";
    tmp(71509) := x"2104";
    tmp(71510) := x"1903";
    tmp(71511) := x"1903";
    tmp(71512) := x"18e3";
    tmp(71513) := x"18e3";
    tmp(71514) := x"18c3";
    tmp(71515) := x"18c2";
    tmp(71516) := x"10c2";
    tmp(71517) := x"10c2";
    tmp(71518) := x"10a2";
    tmp(71519) := x"10a2";
    tmp(71520) := x"0000";
    tmp(71521) := x"0021";
    tmp(71522) := x"0021";
    tmp(71523) := x"0021";
    tmp(71524) := x"0021";
    tmp(71525) := x"0021";
    tmp(71526) := x"0041";
    tmp(71527) := x"0041";
    tmp(71528) := x"0041";
    tmp(71529) := x"0041";
    tmp(71530) := x"0041";
    tmp(71531) := x"0041";
    tmp(71532) := x"0061";
    tmp(71533) := x"0041";
    tmp(71534) := x"0041";
    tmp(71535) := x"0041";
    tmp(71536) := x"0041";
    tmp(71537) := x"0041";
    tmp(71538) := x"0041";
    tmp(71539) := x"0041";
    tmp(71540) := x"0041";
    tmp(71541) := x"0041";
    tmp(71542) := x"0021";
    tmp(71543) := x"0020";
    tmp(71544) := x"0020";
    tmp(71545) := x"0020";
    tmp(71546) := x"0041";
    tmp(71547) := x"0041";
    tmp(71548) := x"0041";
    tmp(71549) := x"0041";
    tmp(71550) := x"0041";
    tmp(71551) := x"0041";
    tmp(71552) := x"0061";
    tmp(71553) := x"0061";
    tmp(71554) := x"0061";
    tmp(71555) := x"0061";
    tmp(71556) := x"0061";
    tmp(71557) := x"0041";
    tmp(71558) := x"0041";
    tmp(71559) := x"0061";
    tmp(71560) := x"0062";
    tmp(71561) := x"0041";
    tmp(71562) := x"0041";
    tmp(71563) := x"0040";
    tmp(71564) := x"0040";
    tmp(71565) := x"0040";
    tmp(71566) := x"0040";
    tmp(71567) := x"0040";
    tmp(71568) := x"0040";
    tmp(71569) := x"0040";
    tmp(71570) := x"0040";
    tmp(71571) := x"0040";
    tmp(71572) := x"0040";
    tmp(71573) := x"0040";
    tmp(71574) := x"0040";
    tmp(71575) := x"0040";
    tmp(71576) := x"0040";
    tmp(71577) := x"0040";
    tmp(71578) := x"0040";
    tmp(71579) := x"0040";
    tmp(71580) := x"0040";
    tmp(71581) := x"0040";
    tmp(71582) := x"0040";
    tmp(71583) := x"0040";
    tmp(71584) := x"0040";
    tmp(71585) := x"0040";
    tmp(71586) := x"0040";
    tmp(71587) := x"0040";
    tmp(71588) := x"0040";
    tmp(71589) := x"0060";
    tmp(71590) := x"0060";
    tmp(71591) := x"0060";
    tmp(71592) := x"0040";
    tmp(71593) := x"0860";
    tmp(71594) := x"0860";
    tmp(71595) := x"0840";
    tmp(71596) := x"0840";
    tmp(71597) := x"0840";
    tmp(71598) := x"0840";
    tmp(71599) := x"0840";
    tmp(71600) := x"0840";
    tmp(71601) := x"0840";
    tmp(71602) := x"0820";
    tmp(71603) := x"0820";
    tmp(71604) := x"0820";
    tmp(71605) := x"0800";
    tmp(71606) := x"1000";
    tmp(71607) := x"1800";
    tmp(71608) := x"1800";
    tmp(71609) := x"1800";
    tmp(71610) := x"2000";
    tmp(71611) := x"1800";
    tmp(71612) := x"2000";
    tmp(71613) := x"2800";
    tmp(71614) := x"2000";
    tmp(71615) := x"2800";
    tmp(71616) := x"2020";
    tmp(71617) := x"2020";
    tmp(71618) := x"1820";
    tmp(71619) := x"1820";
    tmp(71620) := x"2000";
    tmp(71621) := x"2000";
    tmp(71622) := x"3020";
    tmp(71623) := x"4020";
    tmp(71624) := x"4020";
    tmp(71625) := x"4840";
    tmp(71626) := x"4020";
    tmp(71627) := x"3020";
    tmp(71628) := x"3820";
    tmp(71629) := x"4020";
    tmp(71630) := x"4820";
    tmp(71631) := x"4820";
    tmp(71632) := x"4020";
    tmp(71633) := x"4000";
    tmp(71634) := x"4820";
    tmp(71635) := x"3000";
    tmp(71636) := x"3800";
    tmp(71637) := x"4020";
    tmp(71638) := x"4020";
    tmp(71639) := x"3820";
    tmp(71640) := x"4020";
    tmp(71641) := x"2000";
    tmp(71642) := x"2800";
    tmp(71643) := x"3800";
    tmp(71644) := x"3000";
    tmp(71645) := x"3000";
    tmp(71646) := x"3000";
    tmp(71647) := x"2800";
    tmp(71648) := x"2000";
    tmp(71649) := x"1800";
    tmp(71650) := x"2041";
    tmp(71651) := x"20a2";
    tmp(71652) := x"20a1";
    tmp(71653) := x"2081";
    tmp(71654) := x"20c2";
    tmp(71655) := x"18c2";
    tmp(71656) := x"18a2";
    tmp(71657) := x"18c2";
    tmp(71658) := x"18c2";
    tmp(71659) := x"18c2";
    tmp(71660) := x"18a2";
    tmp(71661) := x"18a2";
    tmp(71662) := x"18a2";
    tmp(71663) := x"18a2";
    tmp(71664) := x"18a1";
    tmp(71665) := x"18a1";
    tmp(71666) := x"18a1";
    tmp(71667) := x"10a1";
    tmp(71668) := x"10a1";
    tmp(71669) := x"1081";
    tmp(71670) := x"1081";
    tmp(71671) := x"1081";
    tmp(71672) := x"1081";
    tmp(71673) := x"1081";
    tmp(71674) := x"1061";
    tmp(71675) := x"1061";
    tmp(71676) := x"1061";
    tmp(71677) := x"1061";
    tmp(71678) := x"1061";
    tmp(71679) := x"0841";
    tmp(71680) := x"0840";
    tmp(71681) := x"0840";
    tmp(71682) := x"0840";
    tmp(71683) := x"0840";
    tmp(71684) := x"0840";
    tmp(71685) := x"0840";
    tmp(71686) := x"0840";
    tmp(71687) := x"0820";
    tmp(71688) := x"0820";
    tmp(71689) := x"0820";
    tmp(71690) := x"0820";
    tmp(71691) := x"0820";
    tmp(71692) := x"0820";
    tmp(71693) := x"0820";
    tmp(71694) := x"0820";
    tmp(71695) := x"0020";
    tmp(71696) := x"0020";
    tmp(71697) := x"0020";
    tmp(71698) := x"0020";
    tmp(71699) := x"0020";
    tmp(71700) := x"0020";
    tmp(71701) := x"0020";
    tmp(71702) := x"0020";
    tmp(71703) := x"0020";
    tmp(71704) := x"0020";
    tmp(71705) := x"0000";
    tmp(71706) := x"0000";
    tmp(71707) := x"0000";
    tmp(71708) := x"0000";
    tmp(71709) := x"0020";
    tmp(71710) := x"0020";
    tmp(71711) := x"0020";
    tmp(71712) := x"0020";
    tmp(71713) := x"0020";
    tmp(71714) := x"0020";
    tmp(71715) := x"0020";
    tmp(71716) := x"0020";
    tmp(71717) := x"0020";
    tmp(71718) := x"0020";
    tmp(71719) := x"0820";
    tmp(71720) := x"0820";
    tmp(71721) := x"0820";
    tmp(71722) := x"0820";
    tmp(71723) := x"0820";
    tmp(71724) := x"0840";
    tmp(71725) := x"0840";
    tmp(71726) := x"0840";
    tmp(71727) := x"0841";
    tmp(71728) := x"0861";
    tmp(71729) := x"0861";
    tmp(71730) := x"1081";
    tmp(71731) := x"1081";
    tmp(71732) := x"1081";
    tmp(71733) := x"10a2";
    tmp(71734) := x"10a2";
    tmp(71735) := x"18c2";
    tmp(71736) := x"18c2";
    tmp(71737) := x"18e3";
    tmp(71738) := x"18c3";
    tmp(71739) := x"18e3";
    tmp(71740) := x"18e3";
    tmp(71741) := x"18e3";
    tmp(71742) := x"18e3";
    tmp(71743) := x"18e3";
    tmp(71744) := x"18e3";
    tmp(71745) := x"18e3";
    tmp(71746) := x"18e3";
    tmp(71747) := x"18e3";
    tmp(71748) := x"18c3";
    tmp(71749) := x"18c3";
    tmp(71750) := x"18c3";
    tmp(71751) := x"18c2";
    tmp(71752) := x"18c2";
    tmp(71753) := x"10a2";
    tmp(71754) := x"10a2";
    tmp(71755) := x"10a2";
    tmp(71756) := x"10a2";
    tmp(71757) := x"10a2";
    tmp(71758) := x"1081";
    tmp(71759) := x"1081";
    tmp(71760) := x"0000";
    tmp(71761) := x"0021";
    tmp(71762) := x"0021";
    tmp(71763) := x"0021";
    tmp(71764) := x"0021";
    tmp(71765) := x"0021";
    tmp(71766) := x"0041";
    tmp(71767) := x"0041";
    tmp(71768) := x"0041";
    tmp(71769) := x"0041";
    tmp(71770) := x"0041";
    tmp(71771) := x"0041";
    tmp(71772) := x"0041";
    tmp(71773) := x"0041";
    tmp(71774) := x"0041";
    tmp(71775) := x"0041";
    tmp(71776) := x"0041";
    tmp(71777) := x"0041";
    tmp(71778) := x"0041";
    tmp(71779) := x"0041";
    tmp(71780) := x"0041";
    tmp(71781) := x"0021";
    tmp(71782) := x"0020";
    tmp(71783) := x"0020";
    tmp(71784) := x"0020";
    tmp(71785) := x"0020";
    tmp(71786) := x"0020";
    tmp(71787) := x"0041";
    tmp(71788) := x"0041";
    tmp(71789) := x"0041";
    tmp(71790) := x"0041";
    tmp(71791) := x"0041";
    tmp(71792) := x"0041";
    tmp(71793) := x"0061";
    tmp(71794) := x"0061";
    tmp(71795) := x"0061";
    tmp(71796) := x"0041";
    tmp(71797) := x"0021";
    tmp(71798) := x"0041";
    tmp(71799) := x"0061";
    tmp(71800) := x"0061";
    tmp(71801) := x"0061";
    tmp(71802) := x"0041";
    tmp(71803) := x"0041";
    tmp(71804) := x"0041";
    tmp(71805) := x"0061";
    tmp(71806) := x"0061";
    tmp(71807) := x"0040";
    tmp(71808) := x"0040";
    tmp(71809) := x"0040";
    tmp(71810) := x"0040";
    tmp(71811) := x"0040";
    tmp(71812) := x"0040";
    tmp(71813) := x"0040";
    tmp(71814) := x"0040";
    tmp(71815) := x"0040";
    tmp(71816) := x"0040";
    tmp(71817) := x"0040";
    tmp(71818) := x"0040";
    tmp(71819) := x"0040";
    tmp(71820) := x"0040";
    tmp(71821) := x"0040";
    tmp(71822) := x"0040";
    tmp(71823) := x"0040";
    tmp(71824) := x"0040";
    tmp(71825) := x"0040";
    tmp(71826) := x"0040";
    tmp(71827) := x"0040";
    tmp(71828) := x"0040";
    tmp(71829) := x"0040";
    tmp(71830) := x"0040";
    tmp(71831) := x"0060";
    tmp(71832) := x"0060";
    tmp(71833) := x"0860";
    tmp(71834) := x"0840";
    tmp(71835) := x"0840";
    tmp(71836) := x"0840";
    tmp(71837) := x"0840";
    tmp(71838) := x"0840";
    tmp(71839) := x"0840";
    tmp(71840) := x"0040";
    tmp(71841) := x"0040";
    tmp(71842) := x"0840";
    tmp(71843) := x"0820";
    tmp(71844) := x"0800";
    tmp(71845) := x"0800";
    tmp(71846) := x"1000";
    tmp(71847) := x"1800";
    tmp(71848) := x"1800";
    tmp(71849) := x"2000";
    tmp(71850) := x"2800";
    tmp(71851) := x"2800";
    tmp(71852) := x"2800";
    tmp(71853) := x"3000";
    tmp(71854) := x"3000";
    tmp(71855) := x"3000";
    tmp(71856) := x"3020";
    tmp(71857) := x"3020";
    tmp(71858) := x"2020";
    tmp(71859) := x"1820";
    tmp(71860) := x"1800";
    tmp(71861) := x"1800";
    tmp(71862) := x"2820";
    tmp(71863) := x"3020";
    tmp(71864) := x"3820";
    tmp(71865) := x"4020";
    tmp(71866) := x"3820";
    tmp(71867) := x"3800";
    tmp(71868) := x"4020";
    tmp(71869) := x"4820";
    tmp(71870) := x"4820";
    tmp(71871) := x"4020";
    tmp(71872) := x"3800";
    tmp(71873) := x"4020";
    tmp(71874) := x"3800";
    tmp(71875) := x"3000";
    tmp(71876) := x"3800";
    tmp(71877) := x"3800";
    tmp(71878) := x"3020";
    tmp(71879) := x"2800";
    tmp(71880) := x"3020";
    tmp(71881) := x"2000";
    tmp(71882) := x"3000";
    tmp(71883) := x"3000";
    tmp(71884) := x"3000";
    tmp(71885) := x"3000";
    tmp(71886) := x"3000";
    tmp(71887) := x"2000";
    tmp(71888) := x"2000";
    tmp(71889) := x"1820";
    tmp(71890) := x"20a1";
    tmp(71891) := x"18c2";
    tmp(71892) := x"20a1";
    tmp(71893) := x"20c2";
    tmp(71894) := x"18c2";
    tmp(71895) := x"18c2";
    tmp(71896) := x"18a2";
    tmp(71897) := x"18c2";
    tmp(71898) := x"18a2";
    tmp(71899) := x"18c2";
    tmp(71900) := x"18a1";
    tmp(71901) := x"18a1";
    tmp(71902) := x"18a1";
    tmp(71903) := x"18a1";
    tmp(71904) := x"18a1";
    tmp(71905) := x"18a1";
    tmp(71906) := x"10a1";
    tmp(71907) := x"1081";
    tmp(71908) := x"1081";
    tmp(71909) := x"1081";
    tmp(71910) := x"1081";
    tmp(71911) := x"1081";
    tmp(71912) := x"1081";
    tmp(71913) := x"1061";
    tmp(71914) := x"1061";
    tmp(71915) := x"1061";
    tmp(71916) := x"1061";
    tmp(71917) := x"1061";
    tmp(71918) := x"0841";
    tmp(71919) := x"0840";
    tmp(71920) := x"0840";
    tmp(71921) := x"0840";
    tmp(71922) := x"0840";
    tmp(71923) := x"0840";
    tmp(71924) := x"0840";
    tmp(71925) := x"0840";
    tmp(71926) := x"0820";
    tmp(71927) := x"0820";
    tmp(71928) := x"0820";
    tmp(71929) := x"0820";
    tmp(71930) := x"0820";
    tmp(71931) := x"0020";
    tmp(71932) := x"0020";
    tmp(71933) := x"0020";
    tmp(71934) := x"0020";
    tmp(71935) := x"0020";
    tmp(71936) := x"0020";
    tmp(71937) := x"0020";
    tmp(71938) := x"0020";
    tmp(71939) := x"0020";
    tmp(71940) := x"0020";
    tmp(71941) := x"0000";
    tmp(71942) := x"0000";
    tmp(71943) := x"0000";
    tmp(71944) := x"0000";
    tmp(71945) := x"0000";
    tmp(71946) := x"0000";
    tmp(71947) := x"0000";
    tmp(71948) := x"0000";
    tmp(71949) := x"0000";
    tmp(71950) := x"0020";
    tmp(71951) := x"0020";
    tmp(71952) := x"0020";
    tmp(71953) := x"0020";
    tmp(71954) := x"0020";
    tmp(71955) := x"0020";
    tmp(71956) := x"0020";
    tmp(71957) := x"0020";
    tmp(71958) := x"0020";
    tmp(71959) := x"0020";
    tmp(71960) := x"0020";
    tmp(71961) := x"0020";
    tmp(71962) := x"0820";
    tmp(71963) := x"0820";
    tmp(71964) := x"0820";
    tmp(71965) := x"0820";
    tmp(71966) := x"0820";
    tmp(71967) := x"0840";
    tmp(71968) := x"0840";
    tmp(71969) := x"0840";
    tmp(71970) := x"0841";
    tmp(71971) := x"0861";
    tmp(71972) := x"0861";
    tmp(71973) := x"0861";
    tmp(71974) := x"1081";
    tmp(71975) := x"1081";
    tmp(71976) := x"1081";
    tmp(71977) := x"1082";
    tmp(71978) := x"1082";
    tmp(71979) := x"10a2";
    tmp(71980) := x"10a2";
    tmp(71981) := x"10a2";
    tmp(71982) := x"10a2";
    tmp(71983) := x"10a2";
    tmp(71984) := x"10a2";
    tmp(71985) := x"10a2";
    tmp(71986) := x"10a2";
    tmp(71987) := x"10a2";
    tmp(71988) := x"10a2";
    tmp(71989) := x"10a2";
    tmp(71990) := x"10a2";
    tmp(71991) := x"10a2";
    tmp(71992) := x"10a2";
    tmp(71993) := x"1082";
    tmp(71994) := x"1082";
    tmp(71995) := x"1081";
    tmp(71996) := x"1081";
    tmp(71997) := x"1081";
    tmp(71998) := x"0861";
    tmp(71999) := x"0861";
    tmp(72000) := x"0000";
    tmp(72001) := x"0021";
    tmp(72002) := x"0021";
    tmp(72003) := x"0041";
    tmp(72004) := x"0041";
    tmp(72005) := x"0041";
    tmp(72006) := x"0041";
    tmp(72007) := x"0041";
    tmp(72008) := x"0041";
    tmp(72009) := x"0041";
    tmp(72010) := x"0041";
    tmp(72011) := x"0041";
    tmp(72012) := x"0041";
    tmp(72013) := x"0041";
    tmp(72014) := x"0041";
    tmp(72015) := x"0041";
    tmp(72016) := x"0041";
    tmp(72017) := x"0041";
    tmp(72018) := x"0041";
    tmp(72019) := x"0041";
    tmp(72020) := x"0041";
    tmp(72021) := x"0041";
    tmp(72022) := x"0041";
    tmp(72023) := x"0021";
    tmp(72024) := x"0020";
    tmp(72025) := x"0020";
    tmp(72026) := x"0020";
    tmp(72027) := x"0020";
    tmp(72028) := x"0040";
    tmp(72029) := x"0040";
    tmp(72030) := x"0041";
    tmp(72031) := x"0041";
    tmp(72032) := x"0041";
    tmp(72033) := x"0041";
    tmp(72034) := x"0041";
    tmp(72035) := x"0041";
    tmp(72036) := x"0020";
    tmp(72037) := x"0021";
    tmp(72038) := x"0041";
    tmp(72039) := x"0041";
    tmp(72040) := x"0061";
    tmp(72041) := x"0061";
    tmp(72042) := x"0061";
    tmp(72043) := x"0061";
    tmp(72044) := x"0041";
    tmp(72045) := x"0061";
    tmp(72046) := x"0061";
    tmp(72047) := x"0061";
    tmp(72048) := x"0040";
    tmp(72049) := x"0040";
    tmp(72050) := x"0040";
    tmp(72051) := x"0060";
    tmp(72052) := x"0060";
    tmp(72053) := x"0060";
    tmp(72054) := x"0060";
    tmp(72055) := x"0060";
    tmp(72056) := x"0040";
    tmp(72057) := x"0040";
    tmp(72058) := x"0040";
    tmp(72059) := x"0040";
    tmp(72060) := x"0040";
    tmp(72061) := x"0040";
    tmp(72062) := x"0040";
    tmp(72063) := x"0040";
    tmp(72064) := x"0040";
    tmp(72065) := x"0040";
    tmp(72066) := x"0040";
    tmp(72067) := x"0040";
    tmp(72068) := x"0040";
    tmp(72069) := x"0040";
    tmp(72070) := x"0060";
    tmp(72071) := x"0060";
    tmp(72072) := x"0040";
    tmp(72073) := x"0040";
    tmp(72074) := x"0040";
    tmp(72075) := x"0840";
    tmp(72076) := x"0840";
    tmp(72077) := x"0840";
    tmp(72078) := x"0840";
    tmp(72079) := x"0840";
    tmp(72080) := x"0840";
    tmp(72081) := x"0840";
    tmp(72082) := x"0820";
    tmp(72083) := x"0820";
    tmp(72084) := x"0800";
    tmp(72085) := x"1000";
    tmp(72086) := x"1800";
    tmp(72087) := x"2000";
    tmp(72088) := x"2800";
    tmp(72089) := x"3020";
    tmp(72090) := x"3020";
    tmp(72091) := x"3020";
    tmp(72092) := x"3020";
    tmp(72093) := x"3020";
    tmp(72094) := x"3820";
    tmp(72095) := x"3020";
    tmp(72096) := x"3020";
    tmp(72097) := x"3020";
    tmp(72098) := x"2800";
    tmp(72099) := x"2800";
    tmp(72100) := x"3020";
    tmp(72101) := x"3020";
    tmp(72102) := x"3020";
    tmp(72103) := x"2800";
    tmp(72104) := x"3000";
    tmp(72105) := x"3000";
    tmp(72106) := x"3000";
    tmp(72107) := x"3800";
    tmp(72108) := x"4020";
    tmp(72109) := x"4820";
    tmp(72110) := x"4820";
    tmp(72111) := x"4020";
    tmp(72112) := x"3820";
    tmp(72113) := x"4020";
    tmp(72114) := x"3000";
    tmp(72115) := x"3000";
    tmp(72116) := x"3000";
    tmp(72117) := x"2820";
    tmp(72118) := x"2820";
    tmp(72119) := x"3020";
    tmp(72120) := x"2820";
    tmp(72121) := x"2800";
    tmp(72122) := x"3000";
    tmp(72123) := x"2800";
    tmp(72124) := x"2800";
    tmp(72125) := x"2800";
    tmp(72126) := x"2000";
    tmp(72127) := x"2000";
    tmp(72128) := x"2041";
    tmp(72129) := x"1881";
    tmp(72130) := x"18a1";
    tmp(72131) := x"18a1";
    tmp(72132) := x"18a2";
    tmp(72133) := x"18c2";
    tmp(72134) := x"18a2";
    tmp(72135) := x"18a2";
    tmp(72136) := x"18a2";
    tmp(72137) := x"18a2";
    tmp(72138) := x"18a1";
    tmp(72139) := x"18a1";
    tmp(72140) := x"18a1";
    tmp(72141) := x"18a1";
    tmp(72142) := x"18a1";
    tmp(72143) := x"18a1";
    tmp(72144) := x"10a1";
    tmp(72145) := x"10a1";
    tmp(72146) := x"10a1";
    tmp(72147) := x"1081";
    tmp(72148) := x"1081";
    tmp(72149) := x"1081";
    tmp(72150) := x"1081";
    tmp(72151) := x"1081";
    tmp(72152) := x"1061";
    tmp(72153) := x"1061";
    tmp(72154) := x"1061";
    tmp(72155) := x"1061";
    tmp(72156) := x"0861";
    tmp(72157) := x"0860";
    tmp(72158) := x"0860";
    tmp(72159) := x"0840";
    tmp(72160) := x"0840";
    tmp(72161) := x"0840";
    tmp(72162) := x"0840";
    tmp(72163) := x"0840";
    tmp(72164) := x"0840";
    tmp(72165) := x"0820";
    tmp(72166) := x"0820";
    tmp(72167) := x"0820";
    tmp(72168) := x"0820";
    tmp(72169) := x"0820";
    tmp(72170) := x"0020";
    tmp(72171) := x"0020";
    tmp(72172) := x"0020";
    tmp(72173) := x"0020";
    tmp(72174) := x"0020";
    tmp(72175) := x"0020";
    tmp(72176) := x"0020";
    tmp(72177) := x"0020";
    tmp(72178) := x"0020";
    tmp(72179) := x"0000";
    tmp(72180) := x"0000";
    tmp(72181) := x"0020";
    tmp(72182) := x"0000";
    tmp(72183) := x"0000";
    tmp(72184) := x"0020";
    tmp(72185) := x"0000";
    tmp(72186) := x"0000";
    tmp(72187) := x"0000";
    tmp(72188) := x"0000";
    tmp(72189) := x"0000";
    tmp(72190) := x"0000";
    tmp(72191) := x"0020";
    tmp(72192) := x"0020";
    tmp(72193) := x"0020";
    tmp(72194) := x"0020";
    tmp(72195) := x"0020";
    tmp(72196) := x"0020";
    tmp(72197) := x"0020";
    tmp(72198) := x"0020";
    tmp(72199) := x"0020";
    tmp(72200) := x"0020";
    tmp(72201) := x"0020";
    tmp(72202) := x"0020";
    tmp(72203) := x"0020";
    tmp(72204) := x"0820";
    tmp(72205) := x"0820";
    tmp(72206) := x"0820";
    tmp(72207) := x"0820";
    tmp(72208) := x"0820";
    tmp(72209) := x"0820";
    tmp(72210) := x"0820";
    tmp(72211) := x"0840";
    tmp(72212) := x"0840";
    tmp(72213) := x"0841";
    tmp(72214) := x"0841";
    tmp(72215) := x"0861";
    tmp(72216) := x"0861";
    tmp(72217) := x"0861";
    tmp(72218) := x"0861";
    tmp(72219) := x"1061";
    tmp(72220) := x"1081";
    tmp(72221) := x"1081";
    tmp(72222) := x"1081";
    tmp(72223) := x"1081";
    tmp(72224) := x"1081";
    tmp(72225) := x"1082";
    tmp(72226) := x"1082";
    tmp(72227) := x"1082";
    tmp(72228) := x"1082";
    tmp(72229) := x"1082";
    tmp(72230) := x"1081";
    tmp(72231) := x"1081";
    tmp(72232) := x"1081";
    tmp(72233) := x"0881";
    tmp(72234) := x"0861";
    tmp(72235) := x"0861";
    tmp(72236) := x"0861";
    tmp(72237) := x"0861";
    tmp(72238) := x"0861";
    tmp(72239) := x"0841";
    tmp(72240) := x"0000";
    tmp(72241) := x"0041";
    tmp(72242) := x"0041";
    tmp(72243) := x"0041";
    tmp(72244) := x"0041";
    tmp(72245) := x"0041";
    tmp(72246) := x"0041";
    tmp(72247) := x"0041";
    tmp(72248) := x"0041";
    tmp(72249) := x"0041";
    tmp(72250) := x"0041";
    tmp(72251) := x"0041";
    tmp(72252) := x"0041";
    tmp(72253) := x"0041";
    tmp(72254) := x"0041";
    tmp(72255) := x"0041";
    tmp(72256) := x"0041";
    tmp(72257) := x"0041";
    tmp(72258) := x"0041";
    tmp(72259) := x"0041";
    tmp(72260) := x"0041";
    tmp(72261) := x"0041";
    tmp(72262) := x"0041";
    tmp(72263) := x"0041";
    tmp(72264) := x"0041";
    tmp(72265) := x"0041";
    tmp(72266) := x"0040";
    tmp(72267) := x"0040";
    tmp(72268) := x"0040";
    tmp(72269) := x"0040";
    tmp(72270) := x"0040";
    tmp(72271) := x"0040";
    tmp(72272) := x"0040";
    tmp(72273) := x"0040";
    tmp(72274) := x"0040";
    tmp(72275) := x"0020";
    tmp(72276) := x"0021";
    tmp(72277) := x"0041";
    tmp(72278) := x"0041";
    tmp(72279) := x"0041";
    tmp(72280) := x"0061";
    tmp(72281) := x"0061";
    tmp(72282) := x"0061";
    tmp(72283) := x"0061";
    tmp(72284) := x"0062";
    tmp(72285) := x"0061";
    tmp(72286) := x"0061";
    tmp(72287) := x"0061";
    tmp(72288) := x"0061";
    tmp(72289) := x"0060";
    tmp(72290) := x"0040";
    tmp(72291) := x"0040";
    tmp(72292) := x"0060";
    tmp(72293) := x"0060";
    tmp(72294) := x"0060";
    tmp(72295) := x"0060";
    tmp(72296) := x"0060";
    tmp(72297) := x"0060";
    tmp(72298) := x"0040";
    tmp(72299) := x"0040";
    tmp(72300) := x"0040";
    tmp(72301) := x"0040";
    tmp(72302) := x"0040";
    tmp(72303) := x"0040";
    tmp(72304) := x"0040";
    tmp(72305) := x"0040";
    tmp(72306) := x"0040";
    tmp(72307) := x"0040";
    tmp(72308) := x"0040";
    tmp(72309) := x"0060";
    tmp(72310) := x"0060";
    tmp(72311) := x"0040";
    tmp(72312) := x"0040";
    tmp(72313) := x"0040";
    tmp(72314) := x"0040";
    tmp(72315) := x"0840";
    tmp(72316) := x"0840";
    tmp(72317) := x"0840";
    tmp(72318) := x"0840";
    tmp(72319) := x"0840";
    tmp(72320) := x"0840";
    tmp(72321) := x"0820";
    tmp(72322) := x"0820";
    tmp(72323) := x"1020";
    tmp(72324) := x"1800";
    tmp(72325) := x"2000";
    tmp(72326) := x"2800";
    tmp(72327) := x"2800";
    tmp(72328) := x"2820";
    tmp(72329) := x"3020";
    tmp(72330) := x"3020";
    tmp(72331) := x"3020";
    tmp(72332) := x"3020";
    tmp(72333) := x"2820";
    tmp(72334) := x"2820";
    tmp(72335) := x"2020";
    tmp(72336) := x"1800";
    tmp(72337) := x"1800";
    tmp(72338) := x"2000";
    tmp(72339) := x"2800";
    tmp(72340) := x"2800";
    tmp(72341) := x"2800";
    tmp(72342) := x"2800";
    tmp(72343) := x"2800";
    tmp(72344) := x"3000";
    tmp(72345) := x"2800";
    tmp(72346) := x"2800";
    tmp(72347) := x"3000";
    tmp(72348) := x"4000";
    tmp(72349) := x"4020";
    tmp(72350) := x"4820";
    tmp(72351) := x"4020";
    tmp(72352) := x"3820";
    tmp(72353) := x"2800";
    tmp(72354) := x"2000";
    tmp(72355) := x"2000";
    tmp(72356) := x"2000";
    tmp(72357) := x"2820";
    tmp(72358) := x"4020";
    tmp(72359) := x"4020";
    tmp(72360) := x"2000";
    tmp(72361) := x"2800";
    tmp(72362) := x"2800";
    tmp(72363) := x"2000";
    tmp(72364) := x"2800";
    tmp(72365) := x"2000";
    tmp(72366) := x"1820";
    tmp(72367) := x"1841";
    tmp(72368) := x"1881";
    tmp(72369) := x"10a1";
    tmp(72370) := x"10a1";
    tmp(72371) := x"10a1";
    tmp(72372) := x"10a1";
    tmp(72373) := x"18a1";
    tmp(72374) := x"18a1";
    tmp(72375) := x"18a1";
    tmp(72376) := x"18a1";
    tmp(72377) := x"18a1";
    tmp(72378) := x"18a1";
    tmp(72379) := x"18a1";
    tmp(72380) := x"18a1";
    tmp(72381) := x"18a1";
    tmp(72382) := x"10a1";
    tmp(72383) := x"10a1";
    tmp(72384) := x"10a1";
    tmp(72385) := x"10a1";
    tmp(72386) := x"1081";
    tmp(72387) := x"1081";
    tmp(72388) := x"1081";
    tmp(72389) := x"1081";
    tmp(72390) := x"1081";
    tmp(72391) := x"1061";
    tmp(72392) := x"1061";
    tmp(72393) := x"1061";
    tmp(72394) := x"1061";
    tmp(72395) := x"1061";
    tmp(72396) := x"0841";
    tmp(72397) := x"0840";
    tmp(72398) := x"0840";
    tmp(72399) := x"0840";
    tmp(72400) := x"0840";
    tmp(72401) := x"0840";
    tmp(72402) := x"0840";
    tmp(72403) := x"0840";
    tmp(72404) := x"0820";
    tmp(72405) := x"0820";
    tmp(72406) := x"0820";
    tmp(72407) := x"0820";
    tmp(72408) := x"0820";
    tmp(72409) := x"0820";
    tmp(72410) := x"0020";
    tmp(72411) := x"0020";
    tmp(72412) := x"0020";
    tmp(72413) := x"0020";
    tmp(72414) := x"0020";
    tmp(72415) := x"0020";
    tmp(72416) := x"0020";
    tmp(72417) := x"0020";
    tmp(72418) := x"0020";
    tmp(72419) := x"0000";
    tmp(72420) := x"0000";
    tmp(72421) := x"0000";
    tmp(72422) := x"0000";
    tmp(72423) := x"0000";
    tmp(72424) := x"0000";
    tmp(72425) := x"0000";
    tmp(72426) := x"0000";
    tmp(72427) := x"0000";
    tmp(72428) := x"0000";
    tmp(72429) := x"0000";
    tmp(72430) := x"0000";
    tmp(72431) := x"0000";
    tmp(72432) := x"0020";
    tmp(72433) := x"0020";
    tmp(72434) := x"0020";
    tmp(72435) := x"0020";
    tmp(72436) := x"0020";
    tmp(72437) := x"0020";
    tmp(72438) := x"0020";
    tmp(72439) := x"0020";
    tmp(72440) := x"0020";
    tmp(72441) := x"0020";
    tmp(72442) := x"0020";
    tmp(72443) := x"0020";
    tmp(72444) := x"0020";
    tmp(72445) := x"0020";
    tmp(72446) := x"0020";
    tmp(72447) := x"0820";
    tmp(72448) := x"0820";
    tmp(72449) := x"0820";
    tmp(72450) := x"0820";
    tmp(72451) := x"0820";
    tmp(72452) := x"0820";
    tmp(72453) := x"0820";
    tmp(72454) := x"0840";
    tmp(72455) := x"0840";
    tmp(72456) := x"0840";
    tmp(72457) := x"0841";
    tmp(72458) := x"0841";
    tmp(72459) := x"0841";
    tmp(72460) := x"0861";
    tmp(72461) := x"0861";
    tmp(72462) := x"0861";
    tmp(72463) := x"0861";
    tmp(72464) := x"0861";
    tmp(72465) := x"0861";
    tmp(72466) := x"0861";
    tmp(72467) := x"0861";
    tmp(72468) := x"0861";
    tmp(72469) := x"0861";
    tmp(72470) := x"0861";
    tmp(72471) := x"0861";
    tmp(72472) := x"0861";
    tmp(72473) := x"0861";
    tmp(72474) := x"0841";
    tmp(72475) := x"0841";
    tmp(72476) := x"0840";
    tmp(72477) := x"0840";
    tmp(72478) := x"0840";
    tmp(72479) := x"0820";
    tmp(72480) := x"0000";
    tmp(72481) := x"0041";
    tmp(72482) := x"0041";
    tmp(72483) := x"0041";
    tmp(72484) := x"0041";
    tmp(72485) := x"0041";
    tmp(72486) := x"0021";
    tmp(72487) := x"0021";
    tmp(72488) := x"0021";
    tmp(72489) := x"0041";
    tmp(72490) := x"0041";
    tmp(72491) := x"0041";
    tmp(72492) := x"0041";
    tmp(72493) := x"0041";
    tmp(72494) := x"0041";
    tmp(72495) := x"0041";
    tmp(72496) := x"0041";
    tmp(72497) := x"0041";
    tmp(72498) := x"0041";
    tmp(72499) := x"0041";
    tmp(72500) := x"0041";
    tmp(72501) := x"0041";
    tmp(72502) := x"0041";
    tmp(72503) := x"0041";
    tmp(72504) := x"0041";
    tmp(72505) := x"0041";
    tmp(72506) := x"0041";
    tmp(72507) := x"0041";
    tmp(72508) := x"0041";
    tmp(72509) := x"0040";
    tmp(72510) := x"0040";
    tmp(72511) := x"0040";
    tmp(72512) := x"0040";
    tmp(72513) := x"0040";
    tmp(72514) := x"0040";
    tmp(72515) := x"0040";
    tmp(72516) := x"0020";
    tmp(72517) := x"0041";
    tmp(72518) := x"0041";
    tmp(72519) := x"0041";
    tmp(72520) := x"0041";
    tmp(72521) := x"0041";
    tmp(72522) := x"0061";
    tmp(72523) := x"0061";
    tmp(72524) := x"0082";
    tmp(72525) := x"0082";
    tmp(72526) := x"0062";
    tmp(72527) := x"0061";
    tmp(72528) := x"0081";
    tmp(72529) := x"0081";
    tmp(72530) := x"0060";
    tmp(72531) := x"0060";
    tmp(72532) := x"0060";
    tmp(72533) := x"0040";
    tmp(72534) := x"0040";
    tmp(72535) := x"0040";
    tmp(72536) := x"0040";
    tmp(72537) := x"0060";
    tmp(72538) := x"0060";
    tmp(72539) := x"0060";
    tmp(72540) := x"0060";
    tmp(72541) := x"0040";
    tmp(72542) := x"0040";
    tmp(72543) := x"0040";
    tmp(72544) := x"0040";
    tmp(72545) := x"0040";
    tmp(72546) := x"0040";
    tmp(72547) := x"0040";
    tmp(72548) := x"0040";
    tmp(72549) := x"0040";
    tmp(72550) := x"0040";
    tmp(72551) := x"0040";
    tmp(72552) := x"0040";
    tmp(72553) := x"0040";
    tmp(72554) := x"0840";
    tmp(72555) := x"0840";
    tmp(72556) := x"0840";
    tmp(72557) := x"0840";
    tmp(72558) := x"0840";
    tmp(72559) := x"0840";
    tmp(72560) := x"0820";
    tmp(72561) := x"0820";
    tmp(72562) := x"1020";
    tmp(72563) := x"1800";
    tmp(72564) := x"2000";
    tmp(72565) := x"2000";
    tmp(72566) := x"2000";
    tmp(72567) := x"2000";
    tmp(72568) := x"2000";
    tmp(72569) := x"2000";
    tmp(72570) := x"2820";
    tmp(72571) := x"2820";
    tmp(72572) := x"3020";
    tmp(72573) := x"3020";
    tmp(72574) := x"2020";
    tmp(72575) := x"1800";
    tmp(72576) := x"1800";
    tmp(72577) := x"1800";
    tmp(72578) := x"2000";
    tmp(72579) := x"2800";
    tmp(72580) := x"2800";
    tmp(72581) := x"2000";
    tmp(72582) := x"2800";
    tmp(72583) := x"2800";
    tmp(72584) := x"2800";
    tmp(72585) := x"2800";
    tmp(72586) := x"3000";
    tmp(72587) := x"3800";
    tmp(72588) := x"4020";
    tmp(72589) := x"4020";
    tmp(72590) := x"4820";
    tmp(72591) := x"4820";
    tmp(72592) := x"3000";
    tmp(72593) := x"1000";
    tmp(72594) := x"1000";
    tmp(72595) := x"1820";
    tmp(72596) := x"2820";
    tmp(72597) := x"3820";
    tmp(72598) := x"4020";
    tmp(72599) := x"4020";
    tmp(72600) := x"2000";
    tmp(72601) := x"2000";
    tmp(72602) := x"1820";
    tmp(72603) := x"2020";
    tmp(72604) := x"1820";
    tmp(72605) := x"1820";
    tmp(72606) := x"1041";
    tmp(72607) := x"1081";
    tmp(72608) := x"1081";
    tmp(72609) := x"1081";
    tmp(72610) := x"1081";
    tmp(72611) := x"1081";
    tmp(72612) := x"10a1";
    tmp(72613) := x"10a1";
    tmp(72614) := x"10a1";
    tmp(72615) := x"10a1";
    tmp(72616) := x"10a1";
    tmp(72617) := x"10a1";
    tmp(72618) := x"10a1";
    tmp(72619) := x"10a1";
    tmp(72620) := x"10a1";
    tmp(72621) := x"10a1";
    tmp(72622) := x"10a1";
    tmp(72623) := x"10a1";
    tmp(72624) := x"1081";
    tmp(72625) := x"1081";
    tmp(72626) := x"1081";
    tmp(72627) := x"1081";
    tmp(72628) := x"1081";
    tmp(72629) := x"1061";
    tmp(72630) := x"1061";
    tmp(72631) := x"1061";
    tmp(72632) := x"1061";
    tmp(72633) := x"1061";
    tmp(72634) := x"0861";
    tmp(72635) := x"0841";
    tmp(72636) := x"0840";
    tmp(72637) := x"0840";
    tmp(72638) := x"0840";
    tmp(72639) := x"0840";
    tmp(72640) := x"0840";
    tmp(72641) := x"0840";
    tmp(72642) := x"0840";
    tmp(72643) := x"0820";
    tmp(72644) := x"0820";
    tmp(72645) := x"0820";
    tmp(72646) := x"0820";
    tmp(72647) := x"0820";
    tmp(72648) := x"0820";
    tmp(72649) := x"0020";
    tmp(72650) := x"0020";
    tmp(72651) := x"0020";
    tmp(72652) := x"0020";
    tmp(72653) := x"0020";
    tmp(72654) := x"0020";
    tmp(72655) := x"0020";
    tmp(72656) := x"0020";
    tmp(72657) := x"0020";
    tmp(72658) := x"0020";
    tmp(72659) := x"0020";
    tmp(72660) := x"0020";
    tmp(72661) := x"0020";
    tmp(72662) := x"0000";
    tmp(72663) := x"0020";
    tmp(72664) := x"0000";
    tmp(72665) := x"0000";
    tmp(72666) := x"0020";
    tmp(72667) := x"0000";
    tmp(72668) := x"0000";
    tmp(72669) := x"0000";
    tmp(72670) := x"0000";
    tmp(72671) := x"0000";
    tmp(72672) := x"0020";
    tmp(72673) := x"0020";
    tmp(72674) := x"0020";
    tmp(72675) := x"0020";
    tmp(72676) := x"0020";
    tmp(72677) := x"0020";
    tmp(72678) := x"0020";
    tmp(72679) := x"0020";
    tmp(72680) := x"0020";
    tmp(72681) := x"0020";
    tmp(72682) := x"0020";
    tmp(72683) := x"0020";
    tmp(72684) := x"0020";
    tmp(72685) := x"0020";
    tmp(72686) := x"0020";
    tmp(72687) := x"0020";
    tmp(72688) := x"0020";
    tmp(72689) := x"0020";
    tmp(72690) := x"0020";
    tmp(72691) := x"0020";
    tmp(72692) := x"0020";
    tmp(72693) := x"0820";
    tmp(72694) := x"0820";
    tmp(72695) := x"0820";
    tmp(72696) := x"0820";
    tmp(72697) := x"0820";
    tmp(72698) := x"0840";
    tmp(72699) := x"0840";
    tmp(72700) := x"0841";
    tmp(72701) := x"0841";
    tmp(72702) := x"0841";
    tmp(72703) := x"0841";
    tmp(72704) := x"0841";
    tmp(72705) := x"0841";
    tmp(72706) := x"0841";
    tmp(72707) := x"0841";
    tmp(72708) := x"0841";
    tmp(72709) := x"0841";
    tmp(72710) := x"0841";
    tmp(72711) := x"0840";
    tmp(72712) := x"0840";
    tmp(72713) := x"0840";
    tmp(72714) := x"0840";
    tmp(72715) := x"0820";
    tmp(72716) := x"0820";
    tmp(72717) := x"0820";
    tmp(72718) := x"0020";
    tmp(72719) := x"0020";
    tmp(72720) := x"0000";
    tmp(72721) := x"0041";
    tmp(72722) := x"0041";
    tmp(72723) := x"0041";
    tmp(72724) := x"0041";
    tmp(72725) := x"0021";
    tmp(72726) := x"0020";
    tmp(72727) := x"0020";
    tmp(72728) := x"0021";
    tmp(72729) := x"0041";
    tmp(72730) := x"0041";
    tmp(72731) := x"0041";
    tmp(72732) := x"0041";
    tmp(72733) := x"0041";
    tmp(72734) := x"0041";
    tmp(72735) := x"0041";
    tmp(72736) := x"0041";
    tmp(72737) := x"0041";
    tmp(72738) := x"0041";
    tmp(72739) := x"0041";
    tmp(72740) := x"0041";
    tmp(72741) := x"0041";
    tmp(72742) := x"0041";
    tmp(72743) := x"0041";
    tmp(72744) := x"0041";
    tmp(72745) := x"0041";
    tmp(72746) := x"0041";
    tmp(72747) := x"0041";
    tmp(72748) := x"0041";
    tmp(72749) := x"0041";
    tmp(72750) := x"0040";
    tmp(72751) := x"0040";
    tmp(72752) := x"0040";
    tmp(72753) := x"0040";
    tmp(72754) := x"0040";
    tmp(72755) := x"0020";
    tmp(72756) := x"0020";
    tmp(72757) := x"0020";
    tmp(72758) := x"0021";
    tmp(72759) := x"0041";
    tmp(72760) := x"0041";
    tmp(72761) := x"0041";
    tmp(72762) := x"0041";
    tmp(72763) := x"0061";
    tmp(72764) := x"0061";
    tmp(72765) := x"0061";
    tmp(72766) := x"0061";
    tmp(72767) := x"0061";
    tmp(72768) := x"0081";
    tmp(72769) := x"0081";
    tmp(72770) := x"0081";
    tmp(72771) := x"0081";
    tmp(72772) := x"0061";
    tmp(72773) := x"0060";
    tmp(72774) := x"0060";
    tmp(72775) := x"0040";
    tmp(72776) := x"0040";
    tmp(72777) := x"0040";
    tmp(72778) := x"0040";
    tmp(72779) := x"0040";
    tmp(72780) := x"0040";
    tmp(72781) := x"0060";
    tmp(72782) := x"0060";
    tmp(72783) := x"0040";
    tmp(72784) := x"0040";
    tmp(72785) := x"0040";
    tmp(72786) := x"0040";
    tmp(72787) := x"0040";
    tmp(72788) := x"0040";
    tmp(72789) := x"0040";
    tmp(72790) := x"0040";
    tmp(72791) := x"0040";
    tmp(72792) := x"0840";
    tmp(72793) := x"0840";
    tmp(72794) := x"0840";
    tmp(72795) := x"0840";
    tmp(72796) := x"0840";
    tmp(72797) := x"0840";
    tmp(72798) := x"0840";
    tmp(72799) := x"0840";
    tmp(72800) := x"0820";
    tmp(72801) := x"1020";
    tmp(72802) := x"1000";
    tmp(72803) := x"1800";
    tmp(72804) := x"1800";
    tmp(72805) := x"2000";
    tmp(72806) := x"2000";
    tmp(72807) := x"2000";
    tmp(72808) := x"2000";
    tmp(72809) := x"2000";
    tmp(72810) := x"2820";
    tmp(72811) := x"3020";
    tmp(72812) := x"3020";
    tmp(72813) := x"3020";
    tmp(72814) := x"2000";
    tmp(72815) := x"1800";
    tmp(72816) := x"2000";
    tmp(72817) := x"2000";
    tmp(72818) := x"2000";
    tmp(72819) := x"2800";
    tmp(72820) := x"2000";
    tmp(72821) := x"2000";
    tmp(72822) := x"2800";
    tmp(72823) := x"2800";
    tmp(72824) := x"2800";
    tmp(72825) := x"3000";
    tmp(72826) := x"3000";
    tmp(72827) := x"3820";
    tmp(72828) := x"4020";
    tmp(72829) := x"4820";
    tmp(72830) := x"4820";
    tmp(72831) := x"3820";
    tmp(72832) := x"1800";
    tmp(72833) := x"1000";
    tmp(72834) := x"1800";
    tmp(72835) := x"2820";
    tmp(72836) := x"3020";
    tmp(72837) := x"3820";
    tmp(72838) := x"3820";
    tmp(72839) := x"2820";
    tmp(72840) := x"1820";
    tmp(72841) := x"1820";
    tmp(72842) := x"1040";
    tmp(72843) := x"1041";
    tmp(72844) := x"1041";
    tmp(72845) := x"1061";
    tmp(72846) := x"1061";
    tmp(72847) := x"1061";
    tmp(72848) := x"1061";
    tmp(72849) := x"1061";
    tmp(72850) := x"1081";
    tmp(72851) := x"1081";
    tmp(72852) := x"1081";
    tmp(72853) := x"1081";
    tmp(72854) := x"1081";
    tmp(72855) := x"1081";
    tmp(72856) := x"1081";
    tmp(72857) := x"1081";
    tmp(72858) := x"1081";
    tmp(72859) := x"1081";
    tmp(72860) := x"1081";
    tmp(72861) := x"1081";
    tmp(72862) := x"1081";
    tmp(72863) := x"1081";
    tmp(72864) := x"1081";
    tmp(72865) := x"1081";
    tmp(72866) := x"1081";
    tmp(72867) := x"1061";
    tmp(72868) := x"1081";
    tmp(72869) := x"1061";
    tmp(72870) := x"1061";
    tmp(72871) := x"1061";
    tmp(72872) := x"0861";
    tmp(72873) := x"0861";
    tmp(72874) := x"0840";
    tmp(72875) := x"0840";
    tmp(72876) := x"0840";
    tmp(72877) := x"0840";
    tmp(72878) := x"0840";
    tmp(72879) := x"0840";
    tmp(72880) := x"0840";
    tmp(72881) := x"0840";
    tmp(72882) := x"0820";
    tmp(72883) := x"0820";
    tmp(72884) := x"0820";
    tmp(72885) := x"0820";
    tmp(72886) := x"0820";
    tmp(72887) := x"0020";
    tmp(72888) := x"0020";
    tmp(72889) := x"0020";
    tmp(72890) := x"0020";
    tmp(72891) := x"0020";
    tmp(72892) := x"0020";
    tmp(72893) := x"0020";
    tmp(72894) := x"0020";
    tmp(72895) := x"0020";
    tmp(72896) := x"0020";
    tmp(72897) := x"0020";
    tmp(72898) := x"0020";
    tmp(72899) := x"0020";
    tmp(72900) := x"0000";
    tmp(72901) := x"0020";
    tmp(72902) := x"0000";
    tmp(72903) := x"0020";
    tmp(72904) := x"0020";
    tmp(72905) := x"0020";
    tmp(72906) := x"0020";
    tmp(72907) := x"0000";
    tmp(72908) := x"0000";
    tmp(72909) := x"0000";
    tmp(72910) := x"0000";
    tmp(72911) := x"0020";
    tmp(72912) := x"0020";
    tmp(72913) := x"0000";
    tmp(72914) := x"0020";
    tmp(72915) := x"0020";
    tmp(72916) := x"0020";
    tmp(72917) := x"0020";
    tmp(72918) := x"0020";
    tmp(72919) := x"0020";
    tmp(72920) := x"0020";
    tmp(72921) := x"0020";
    tmp(72922) := x"0020";
    tmp(72923) := x"0020";
    tmp(72924) := x"0020";
    tmp(72925) := x"0020";
    tmp(72926) := x"0020";
    tmp(72927) := x"0020";
    tmp(72928) := x"0020";
    tmp(72929) := x"0020";
    tmp(72930) := x"0020";
    tmp(72931) := x"0020";
    tmp(72932) := x"0020";
    tmp(72933) := x"0020";
    tmp(72934) := x"0020";
    tmp(72935) := x"0020";
    tmp(72936) := x"0820";
    tmp(72937) := x"0820";
    tmp(72938) := x"0820";
    tmp(72939) := x"0820";
    tmp(72940) := x"0820";
    tmp(72941) := x"0820";
    tmp(72942) := x"0820";
    tmp(72943) := x"0820";
    tmp(72944) := x"0840";
    tmp(72945) := x"0840";
    tmp(72946) := x"0840";
    tmp(72947) := x"0840";
    tmp(72948) := x"0820";
    tmp(72949) := x"0820";
    tmp(72950) := x"0820";
    tmp(72951) := x"0820";
    tmp(72952) := x"0820";
    tmp(72953) := x"0820";
    tmp(72954) := x"0820";
    tmp(72955) := x"0020";
    tmp(72956) := x"0020";
    tmp(72957) := x"0020";
    tmp(72958) := x"0020";
    tmp(72959) := x"0020";
    tmp(72960) := x"0000";
    tmp(72961) := x"0041";
    tmp(72962) := x"0041";
    tmp(72963) := x"0041";
    tmp(72964) := x"0021";
    tmp(72965) := x"0020";
    tmp(72966) := x"0020";
    tmp(72967) := x"0021";
    tmp(72968) := x"0021";
    tmp(72969) := x"0041";
    tmp(72970) := x"0041";
    tmp(72971) := x"0041";
    tmp(72972) := x"0041";
    tmp(72973) := x"0041";
    tmp(72974) := x"0041";
    tmp(72975) := x"0041";
    tmp(72976) := x"0041";
    tmp(72977) := x"0041";
    tmp(72978) := x"0041";
    tmp(72979) := x"0041";
    tmp(72980) := x"0041";
    tmp(72981) := x"0041";
    tmp(72982) := x"0041";
    tmp(72983) := x"0041";
    tmp(72984) := x"0041";
    tmp(72985) := x"0041";
    tmp(72986) := x"0061";
    tmp(72987) := x"0061";
    tmp(72988) := x"0041";
    tmp(72989) := x"0041";
    tmp(72990) := x"0041";
    tmp(72991) := x"0041";
    tmp(72992) := x"0040";
    tmp(72993) := x"0040";
    tmp(72994) := x"0020";
    tmp(72995) := x"0020";
    tmp(72996) := x"0020";
    tmp(72997) := x"0020";
    tmp(72998) := x"0020";
    tmp(72999) := x"0040";
    tmp(73000) := x"0041";
    tmp(73001) := x"0041";
    tmp(73002) := x"0041";
    tmp(73003) := x"0041";
    tmp(73004) := x"0041";
    tmp(73005) := x"0061";
    tmp(73006) := x"0061";
    tmp(73007) := x"0061";
    tmp(73008) := x"0061";
    tmp(73009) := x"0061";
    tmp(73010) := x"0061";
    tmp(73011) := x"0061";
    tmp(73012) := x"0081";
    tmp(73013) := x"0081";
    tmp(73014) := x"0881";
    tmp(73015) := x"0060";
    tmp(73016) := x"0060";
    tmp(73017) := x"0040";
    tmp(73018) := x"0040";
    tmp(73019) := x"0040";
    tmp(73020) := x"0040";
    tmp(73021) := x"0040";
    tmp(73022) := x"0040";
    tmp(73023) := x"0040";
    tmp(73024) := x"0020";
    tmp(73025) := x"0040";
    tmp(73026) := x"0040";
    tmp(73027) := x"0040";
    tmp(73028) := x"0040";
    tmp(73029) := x"0840";
    tmp(73030) := x"0860";
    tmp(73031) := x"0840";
    tmp(73032) := x"0840";
    tmp(73033) := x"0840";
    tmp(73034) := x"0840";
    tmp(73035) := x"0840";
    tmp(73036) := x"0840";
    tmp(73037) := x"0840";
    tmp(73038) := x"0840";
    tmp(73039) := x"0840";
    tmp(73040) := x"0820";
    tmp(73041) := x"1020";
    tmp(73042) := x"1800";
    tmp(73043) := x"1800";
    tmp(73044) := x"1800";
    tmp(73045) := x"1800";
    tmp(73046) := x"1800";
    tmp(73047) := x"2000";
    tmp(73048) := x"2820";
    tmp(73049) := x"2820";
    tmp(73050) := x"3020";
    tmp(73051) := x"3820";
    tmp(73052) := x"3020";
    tmp(73053) := x"3020";
    tmp(73054) := x"2000";
    tmp(73055) := x"2000";
    tmp(73056) := x"2000";
    tmp(73057) := x"2000";
    tmp(73058) := x"2000";
    tmp(73059) := x"1800";
    tmp(73060) := x"2000";
    tmp(73061) := x"2800";
    tmp(73062) := x"2800";
    tmp(73063) := x"3000";
    tmp(73064) := x"3000";
    tmp(73065) := x"3820";
    tmp(73066) := x"3820";
    tmp(73067) := x"3820";
    tmp(73068) := x"3820";
    tmp(73069) := x"3820";
    tmp(73070) := x"3820";
    tmp(73071) := x"1800";
    tmp(73072) := x"0800";
    tmp(73073) := x"1000";
    tmp(73074) := x"2000";
    tmp(73075) := x"2800";
    tmp(73076) := x"2800";
    tmp(73077) := x"3020";
    tmp(73078) := x"3020";
    tmp(73079) := x"1820";
    tmp(73080) := x"1020";
    tmp(73081) := x"0840";
    tmp(73082) := x"0840";
    tmp(73083) := x"0841";
    tmp(73084) := x"0841";
    tmp(73085) := x"0841";
    tmp(73086) := x"0841";
    tmp(73087) := x"0841";
    tmp(73088) := x"0861";
    tmp(73089) := x"1061";
    tmp(73090) := x"1061";
    tmp(73091) := x"1061";
    tmp(73092) := x"1061";
    tmp(73093) := x"1061";
    tmp(73094) := x"1061";
    tmp(73095) := x"1081";
    tmp(73096) := x"1081";
    tmp(73097) := x"1081";
    tmp(73098) := x"1081";
    tmp(73099) := x"1081";
    tmp(73100) := x"1081";
    tmp(73101) := x"1081";
    tmp(73102) := x"1081";
    tmp(73103) := x"1081";
    tmp(73104) := x"1081";
    tmp(73105) := x"1081";
    tmp(73106) := x"1061";
    tmp(73107) := x"1061";
    tmp(73108) := x"1061";
    tmp(73109) := x"1061";
    tmp(73110) := x"0861";
    tmp(73111) := x"0861";
    tmp(73112) := x"0860";
    tmp(73113) := x"0840";
    tmp(73114) := x"0840";
    tmp(73115) := x"0840";
    tmp(73116) := x"0840";
    tmp(73117) := x"0840";
    tmp(73118) := x"0840";
    tmp(73119) := x"0840";
    tmp(73120) := x"0820";
    tmp(73121) := x"0820";
    tmp(73122) := x"0820";
    tmp(73123) := x"0820";
    tmp(73124) := x"0820";
    tmp(73125) := x"0820";
    tmp(73126) := x"0820";
    tmp(73127) := x"0020";
    tmp(73128) := x"0020";
    tmp(73129) := x"0020";
    tmp(73130) := x"0020";
    tmp(73131) := x"0020";
    tmp(73132) := x"0020";
    tmp(73133) := x"0020";
    tmp(73134) := x"0020";
    tmp(73135) := x"0020";
    tmp(73136) := x"0020";
    tmp(73137) := x"0020";
    tmp(73138) := x"0000";
    tmp(73139) := x"0020";
    tmp(73140) := x"0000";
    tmp(73141) := x"0000";
    tmp(73142) := x"0020";
    tmp(73143) := x"0020";
    tmp(73144) := x"0000";
    tmp(73145) := x"0000";
    tmp(73146) := x"0000";
    tmp(73147) := x"0020";
    tmp(73148) := x"0000";
    tmp(73149) := x"0000";
    tmp(73150) := x"0000";
    tmp(73151) := x"0000";
    tmp(73152) := x"0000";
    tmp(73153) := x"0020";
    tmp(73154) := x"0000";
    tmp(73155) := x"0020";
    tmp(73156) := x"0020";
    tmp(73157) := x"0020";
    tmp(73158) := x"0020";
    tmp(73159) := x"0020";
    tmp(73160) := x"0020";
    tmp(73161) := x"0020";
    tmp(73162) := x"0020";
    tmp(73163) := x"0020";
    tmp(73164) := x"0020";
    tmp(73165) := x"0020";
    tmp(73166) := x"0020";
    tmp(73167) := x"0020";
    tmp(73168) := x"0020";
    tmp(73169) := x"0020";
    tmp(73170) := x"0020";
    tmp(73171) := x"0020";
    tmp(73172) := x"0020";
    tmp(73173) := x"0020";
    tmp(73174) := x"0020";
    tmp(73175) := x"0020";
    tmp(73176) := x"0020";
    tmp(73177) := x"0020";
    tmp(73178) := x"0020";
    tmp(73179) := x"0020";
    tmp(73180) := x"0020";
    tmp(73181) := x"0020";
    tmp(73182) := x"0020";
    tmp(73183) := x"0020";
    tmp(73184) := x"0020";
    tmp(73185) := x"0020";
    tmp(73186) := x"0020";
    tmp(73187) := x"0020";
    tmp(73188) := x"0020";
    tmp(73189) := x"0020";
    tmp(73190) := x"0020";
    tmp(73191) := x"0020";
    tmp(73192) := x"0020";
    tmp(73193) := x"0020";
    tmp(73194) := x"0020";
    tmp(73195) := x"0020";
    tmp(73196) := x"0020";
    tmp(73197) := x"0000";
    tmp(73198) := x"0000";
    tmp(73199) := x"0020";
    tmp(73200) := x"0000";
    tmp(73201) := x"0041";
    tmp(73202) := x"0041";
    tmp(73203) := x"0041";
    tmp(73204) := x"0021";
    tmp(73205) := x"0020";
    tmp(73206) := x"0020";
    tmp(73207) := x"0021";
    tmp(73208) := x"0021";
    tmp(73209) := x"0041";
    tmp(73210) := x"0041";
    tmp(73211) := x"0041";
    tmp(73212) := x"0041";
    tmp(73213) := x"0041";
    tmp(73214) := x"0041";
    tmp(73215) := x"0041";
    tmp(73216) := x"0041";
    tmp(73217) := x"0041";
    tmp(73218) := x"0041";
    tmp(73219) := x"0041";
    tmp(73220) := x"0041";
    tmp(73221) := x"0041";
    tmp(73222) := x"0041";
    tmp(73223) := x"0041";
    tmp(73224) := x"0041";
    tmp(73225) := x"0041";
    tmp(73226) := x"0061";
    tmp(73227) := x"0041";
    tmp(73228) := x"0041";
    tmp(73229) := x"0061";
    tmp(73230) := x"0041";
    tmp(73231) := x"0040";
    tmp(73232) := x"0040";
    tmp(73233) := x"0040";
    tmp(73234) := x"0020";
    tmp(73235) := x"0020";
    tmp(73236) := x"0020";
    tmp(73237) := x"0040";
    tmp(73238) := x"0040";
    tmp(73239) := x"0040";
    tmp(73240) := x"0040";
    tmp(73241) := x"0040";
    tmp(73242) := x"0040";
    tmp(73243) := x"0040";
    tmp(73244) := x"0041";
    tmp(73245) := x"0041";
    tmp(73246) := x"0041";
    tmp(73247) := x"0041";
    tmp(73248) := x"0041";
    tmp(73249) := x"0041";
    tmp(73250) := x"0041";
    tmp(73251) := x"0041";
    tmp(73252) := x"0041";
    tmp(73253) := x"0041";
    tmp(73254) := x"0041";
    tmp(73255) := x"0041";
    tmp(73256) := x"0061";
    tmp(73257) := x"0060";
    tmp(73258) := x"0060";
    tmp(73259) := x"0040";
    tmp(73260) := x"0040";
    tmp(73261) := x"0040";
    tmp(73262) := x"0040";
    tmp(73263) := x"0040";
    tmp(73264) := x"0040";
    tmp(73265) := x"0040";
    tmp(73266) := x"0040";
    tmp(73267) := x"0040";
    tmp(73268) := x"0860";
    tmp(73269) := x"0860";
    tmp(73270) := x"0840";
    tmp(73271) := x"0840";
    tmp(73272) := x"0840";
    tmp(73273) := x"0840";
    tmp(73274) := x"0840";
    tmp(73275) := x"0040";
    tmp(73276) := x"0040";
    tmp(73277) := x"0040";
    tmp(73278) := x"0040";
    tmp(73279) := x"0840";
    tmp(73280) := x"0820";
    tmp(73281) := x"1020";
    tmp(73282) := x"1000";
    tmp(73283) := x"1000";
    tmp(73284) := x"1000";
    tmp(73285) := x"1820";
    tmp(73286) := x"2020";
    tmp(73287) := x"2820";
    tmp(73288) := x"2820";
    tmp(73289) := x"2820";
    tmp(73290) := x"3020";
    tmp(73291) := x"2820";
    tmp(73292) := x"2820";
    tmp(73293) := x"2000";
    tmp(73294) := x"1800";
    tmp(73295) := x"2000";
    tmp(73296) := x"2000";
    tmp(73297) := x"2000";
    tmp(73298) := x"2000";
    tmp(73299) := x"2000";
    tmp(73300) := x"2800";
    tmp(73301) := x"3000";
    tmp(73302) := x"3820";
    tmp(73303) := x"4020";
    tmp(73304) := x"4820";
    tmp(73305) := x"4020";
    tmp(73306) := x"4820";
    tmp(73307) := x"4020";
    tmp(73308) := x"3820";
    tmp(73309) := x"3820";
    tmp(73310) := x"2820";
    tmp(73311) := x"1000";
    tmp(73312) := x"0800";
    tmp(73313) := x"2000";
    tmp(73314) := x"2800";
    tmp(73315) := x"2800";
    tmp(73316) := x"2820";
    tmp(73317) := x"3020";
    tmp(73318) := x"1820";
    tmp(73319) := x"0820";
    tmp(73320) := x"0820";
    tmp(73321) := x"0820";
    tmp(73322) := x"0840";
    tmp(73323) := x"0840";
    tmp(73324) := x"0840";
    tmp(73325) := x"0840";
    tmp(73326) := x"0840";
    tmp(73327) := x"0840";
    tmp(73328) := x"0841";
    tmp(73329) := x"0861";
    tmp(73330) := x"0861";
    tmp(73331) := x"0861";
    tmp(73332) := x"0861";
    tmp(73333) := x"0861";
    tmp(73334) := x"0861";
    tmp(73335) := x"1061";
    tmp(73336) := x"1061";
    tmp(73337) := x"1061";
    tmp(73338) := x"1061";
    tmp(73339) := x"1061";
    tmp(73340) := x"1061";
    tmp(73341) := x"1061";
    tmp(73342) := x"1061";
    tmp(73343) := x"1061";
    tmp(73344) := x"1061";
    tmp(73345) := x"1061";
    tmp(73346) := x"1061";
    tmp(73347) := x"0861";
    tmp(73348) := x"0861";
    tmp(73349) := x"0861";
    tmp(73350) := x"0861";
    tmp(73351) := x"0860";
    tmp(73352) := x"0840";
    tmp(73353) := x"0840";
    tmp(73354) := x"0840";
    tmp(73355) := x"0840";
    tmp(73356) := x"0840";
    tmp(73357) := x"0840";
    tmp(73358) := x"0840";
    tmp(73359) := x"0820";
    tmp(73360) := x"0820";
    tmp(73361) := x"0820";
    tmp(73362) := x"0820";
    tmp(73363) := x"0820";
    tmp(73364) := x"0820";
    tmp(73365) := x"0820";
    tmp(73366) := x"0020";
    tmp(73367) := x"0020";
    tmp(73368) := x"0020";
    tmp(73369) := x"0020";
    tmp(73370) := x"0020";
    tmp(73371) := x"0020";
    tmp(73372) := x"0020";
    tmp(73373) := x"0020";
    tmp(73374) := x"0020";
    tmp(73375) := x"0020";
    tmp(73376) := x"0000";
    tmp(73377) := x"0000";
    tmp(73378) := x"0020";
    tmp(73379) := x"0000";
    tmp(73380) := x"0000";
    tmp(73381) := x"0000";
    tmp(73382) := x"0000";
    tmp(73383) := x"0000";
    tmp(73384) := x"0000";
    tmp(73385) := x"0020";
    tmp(73386) := x"0000";
    tmp(73387) := x"0020";
    tmp(73388) := x"0000";
    tmp(73389) := x"0000";
    tmp(73390) := x"0000";
    tmp(73391) := x"0000";
    tmp(73392) := x"0020";
    tmp(73393) := x"0000";
    tmp(73394) := x"0000";
    tmp(73395) := x"0000";
    tmp(73396) := x"0000";
    tmp(73397) := x"0020";
    tmp(73398) := x"0020";
    tmp(73399) := x"0020";
    tmp(73400) := x"0020";
    tmp(73401) := x"0020";
    tmp(73402) := x"0020";
    tmp(73403) := x"0020";
    tmp(73404) := x"0020";
    tmp(73405) := x"0020";
    tmp(73406) := x"0020";
    tmp(73407) := x"0020";
    tmp(73408) := x"0020";
    tmp(73409) := x"0020";
    tmp(73410) := x"0020";
    tmp(73411) := x"0020";
    tmp(73412) := x"0020";
    tmp(73413) := x"0020";
    tmp(73414) := x"0020";
    tmp(73415) := x"0020";
    tmp(73416) := x"0020";
    tmp(73417) := x"0020";
    tmp(73418) := x"0020";
    tmp(73419) := x"0020";
    tmp(73420) := x"0020";
    tmp(73421) := x"0020";
    tmp(73422) := x"0020";
    tmp(73423) := x"0020";
    tmp(73424) := x"0020";
    tmp(73425) := x"0020";
    tmp(73426) := x"0020";
    tmp(73427) := x"0020";
    tmp(73428) := x"0000";
    tmp(73429) := x"0000";
    tmp(73430) := x"0000";
    tmp(73431) := x"0000";
    tmp(73432) := x"0000";
    tmp(73433) := x"0000";
    tmp(73434) := x"0000";
    tmp(73435) := x"0000";
    tmp(73436) := x"0000";
    tmp(73437) := x"0000";
    tmp(73438) := x"0000";
    tmp(73439) := x"0000";
    tmp(73440) := x"0000";
    tmp(73441) := x"0041";
    tmp(73442) := x"0041";
    tmp(73443) := x"0041";
    tmp(73444) := x"0021";
    tmp(73445) := x"0020";
    tmp(73446) := x"0020";
    tmp(73447) := x"0020";
    tmp(73448) := x"0020";
    tmp(73449) := x"0021";
    tmp(73450) := x"0021";
    tmp(73451) := x"0021";
    tmp(73452) := x"0041";
    tmp(73453) := x"0041";
    tmp(73454) := x"0041";
    tmp(73455) := x"0061";
    tmp(73456) := x"0041";
    tmp(73457) := x"0061";
    tmp(73458) := x"0061";
    tmp(73459) := x"0041";
    tmp(73460) := x"0061";
    tmp(73461) := x"0061";
    tmp(73462) := x"0061";
    tmp(73463) := x"0061";
    tmp(73464) := x"0061";
    tmp(73465) := x"0061";
    tmp(73466) := x"0061";
    tmp(73467) := x"0061";
    tmp(73468) := x"0061";
    tmp(73469) := x"0061";
    tmp(73470) := x"0061";
    tmp(73471) := x"0061";
    tmp(73472) := x"0040";
    tmp(73473) := x"0040";
    tmp(73474) := x"0040";
    tmp(73475) := x"0020";
    tmp(73476) := x"0020";
    tmp(73477) := x"0040";
    tmp(73478) := x"0040";
    tmp(73479) := x"0040";
    tmp(73480) := x"0041";
    tmp(73481) := x"0040";
    tmp(73482) := x"0040";
    tmp(73483) := x"0040";
    tmp(73484) := x"0040";
    tmp(73485) := x"0040";
    tmp(73486) := x"0041";
    tmp(73487) := x"0041";
    tmp(73488) := x"0041";
    tmp(73489) := x"0041";
    tmp(73490) := x"0041";
    tmp(73491) := x"0041";
    tmp(73492) := x"0041";
    tmp(73493) := x"0041";
    tmp(73494) := x"0041";
    tmp(73495) := x"0041";
    tmp(73496) := x"0040";
    tmp(73497) := x"0020";
    tmp(73498) := x"0020";
    tmp(73499) := x"0020";
    tmp(73500) := x"0040";
    tmp(73501) := x"0040";
    tmp(73502) := x"0040";
    tmp(73503) := x"0040";
    tmp(73504) := x"0040";
    tmp(73505) := x"0040";
    tmp(73506) := x"0040";
    tmp(73507) := x"0040";
    tmp(73508) := x"0040";
    tmp(73509) := x"0040";
    tmp(73510) := x"0040";
    tmp(73511) := x"0040";
    tmp(73512) := x"0040";
    tmp(73513) := x"0040";
    tmp(73514) := x"0040";
    tmp(73515) := x"0040";
    tmp(73516) := x"0040";
    tmp(73517) := x"0040";
    tmp(73518) := x"0040";
    tmp(73519) := x"0040";
    tmp(73520) := x"0820";
    tmp(73521) := x"1020";
    tmp(73522) := x"1000";
    tmp(73523) := x"1000";
    tmp(73524) := x"1820";
    tmp(73525) := x"1820";
    tmp(73526) := x"2020";
    tmp(73527) := x"2020";
    tmp(73528) := x"2020";
    tmp(73529) := x"2820";
    tmp(73530) := x"2820";
    tmp(73531) := x"2820";
    tmp(73532) := x"2020";
    tmp(73533) := x"1800";
    tmp(73534) := x"1800";
    tmp(73535) := x"1800";
    tmp(73536) := x"1800";
    tmp(73537) := x"2000";
    tmp(73538) := x"2000";
    tmp(73539) := x"2800";
    tmp(73540) := x"3020";
    tmp(73541) := x"3820";
    tmp(73542) := x"4020";
    tmp(73543) := x"4020";
    tmp(73544) := x"4020";
    tmp(73545) := x"3820";
    tmp(73546) := x"3820";
    tmp(73547) := x"4820";
    tmp(73548) := x"4020";
    tmp(73549) := x"3020";
    tmp(73550) := x"1800";
    tmp(73551) := x"1000";
    tmp(73552) := x"1800";
    tmp(73553) := x"2800";
    tmp(73554) := x"2800";
    tmp(73555) := x"3020";
    tmp(73556) := x"2820";
    tmp(73557) := x"1820";
    tmp(73558) := x"0820";
    tmp(73559) := x"0820";
    tmp(73560) := x"0820";
    tmp(73561) := x"0820";
    tmp(73562) := x"0820";
    tmp(73563) := x"0820";
    tmp(73564) := x"0820";
    tmp(73565) := x"0820";
    tmp(73566) := x"0840";
    tmp(73567) := x"0840";
    tmp(73568) := x"0840";
    tmp(73569) := x"0840";
    tmp(73570) := x"0840";
    tmp(73571) := x"0840";
    tmp(73572) := x"0840";
    tmp(73573) := x"0861";
    tmp(73574) := x"0861";
    tmp(73575) := x"0861";
    tmp(73576) := x"0861";
    tmp(73577) := x"0861";
    tmp(73578) := x"0861";
    tmp(73579) := x"0861";
    tmp(73580) := x"0861";
    tmp(73581) := x"0861";
    tmp(73582) := x"0861";
    tmp(73583) := x"0861";
    tmp(73584) := x"0861";
    tmp(73585) := x"0861";
    tmp(73586) := x"0841";
    tmp(73587) := x"0841";
    tmp(73588) := x"0841";
    tmp(73589) := x"0840";
    tmp(73590) := x"0840";
    tmp(73591) := x"0840";
    tmp(73592) := x"0840";
    tmp(73593) := x"0840";
    tmp(73594) := x"0840";
    tmp(73595) := x"0840";
    tmp(73596) := x"0840";
    tmp(73597) := x"0840";
    tmp(73598) := x"0820";
    tmp(73599) := x"0820";
    tmp(73600) := x"0820";
    tmp(73601) := x"0820";
    tmp(73602) := x"0820";
    tmp(73603) := x"0820";
    tmp(73604) := x"0020";
    tmp(73605) := x"0020";
    tmp(73606) := x"0020";
    tmp(73607) := x"0020";
    tmp(73608) := x"0020";
    tmp(73609) := x"0020";
    tmp(73610) := x"0020";
    tmp(73611) := x"0020";
    tmp(73612) := x"0000";
    tmp(73613) := x"0020";
    tmp(73614) := x"0020";
    tmp(73615) := x"0020";
    tmp(73616) := x"0000";
    tmp(73617) := x"0000";
    tmp(73618) := x"0000";
    tmp(73619) := x"0000";
    tmp(73620) := x"0020";
    tmp(73621) := x"0000";
    tmp(73622) := x"0020";
    tmp(73623) := x"0000";
    tmp(73624) := x"0000";
    tmp(73625) := x"0000";
    tmp(73626) := x"0000";
    tmp(73627) := x"0020";
    tmp(73628) := x"0000";
    tmp(73629) := x"0000";
    tmp(73630) := x"0000";
    tmp(73631) := x"0000";
    tmp(73632) := x"0000";
    tmp(73633) := x"0000";
    tmp(73634) := x"0000";
    tmp(73635) := x"0000";
    tmp(73636) := x"0020";
    tmp(73637) := x"0000";
    tmp(73638) := x"0020";
    tmp(73639) := x"0020";
    tmp(73640) := x"0020";
    tmp(73641) := x"0020";
    tmp(73642) := x"0020";
    tmp(73643) := x"0020";
    tmp(73644) := x"0020";
    tmp(73645) := x"0020";
    tmp(73646) := x"0020";
    tmp(73647) := x"0020";
    tmp(73648) := x"0020";
    tmp(73649) := x"0020";
    tmp(73650) := x"0020";
    tmp(73651) := x"0020";
    tmp(73652) := x"0020";
    tmp(73653) := x"0020";
    tmp(73654) := x"0020";
    tmp(73655) := x"0020";
    tmp(73656) := x"0020";
    tmp(73657) := x"0020";
    tmp(73658) := x"0020";
    tmp(73659) := x"0020";
    tmp(73660) := x"0020";
    tmp(73661) := x"0020";
    tmp(73662) := x"0000";
    tmp(73663) := x"0000";
    tmp(73664) := x"0000";
    tmp(73665) := x"0000";
    tmp(73666) := x"0000";
    tmp(73667) := x"0000";
    tmp(73668) := x"0000";
    tmp(73669) := x"0000";
    tmp(73670) := x"0000";
    tmp(73671) := x"0000";
    tmp(73672) := x"0000";
    tmp(73673) := x"0000";
    tmp(73674) := x"0000";
    tmp(73675) := x"0000";
    tmp(73676) := x"0000";
    tmp(73677) := x"0000";
    tmp(73678) := x"0000";
    tmp(73679) := x"0000";
    tmp(73680) := x"0000";
    tmp(73681) := x"0020";
    tmp(73682) := x"0020";
    tmp(73683) := x"0020";
    tmp(73684) := x"0021";
    tmp(73685) := x"0020";
    tmp(73686) := x"0020";
    tmp(73687) := x"0020";
    tmp(73688) := x"0020";
    tmp(73689) := x"0020";
    tmp(73690) := x"0020";
    tmp(73691) := x"0021";
    tmp(73692) := x"0021";
    tmp(73693) := x"0021";
    tmp(73694) := x"0021";
    tmp(73695) := x"0041";
    tmp(73696) := x"0041";
    tmp(73697) := x"0041";
    tmp(73698) := x"0061";
    tmp(73699) := x"0061";
    tmp(73700) := x"0061";
    tmp(73701) := x"0061";
    tmp(73702) := x"0061";
    tmp(73703) := x"0061";
    tmp(73704) := x"0061";
    tmp(73705) := x"0061";
    tmp(73706) := x"0061";
    tmp(73707) := x"0061";
    tmp(73708) := x"0061";
    tmp(73709) := x"0061";
    tmp(73710) := x"0061";
    tmp(73711) := x"0061";
    tmp(73712) := x"0061";
    tmp(73713) := x"0040";
    tmp(73714) := x"0040";
    tmp(73715) := x"0040";
    tmp(73716) := x"0040";
    tmp(73717) := x"0040";
    tmp(73718) := x"0040";
    tmp(73719) := x"0041";
    tmp(73720) := x"0041";
    tmp(73721) := x"0040";
    tmp(73722) := x"0040";
    tmp(73723) := x"0040";
    tmp(73724) := x"0040";
    tmp(73725) := x"0040";
    tmp(73726) := x"0040";
    tmp(73727) := x"0041";
    tmp(73728) := x"0041";
    tmp(73729) := x"0040";
    tmp(73730) := x"0040";
    tmp(73731) := x"0041";
    tmp(73732) := x"0040";
    tmp(73733) := x"0020";
    tmp(73734) := x"0020";
    tmp(73735) := x"0020";
    tmp(73736) := x"0040";
    tmp(73737) := x"0040";
    tmp(73738) := x"0040";
    tmp(73739) := x"0040";
    tmp(73740) := x"0040";
    tmp(73741) := x"0040";
    tmp(73742) := x"0040";
    tmp(73743) := x"0040";
    tmp(73744) := x"0040";
    tmp(73745) := x"0040";
    tmp(73746) := x"0020";
    tmp(73747) := x"0040";
    tmp(73748) := x"0040";
    tmp(73749) := x"0040";
    tmp(73750) := x"0040";
    tmp(73751) := x"0040";
    tmp(73752) := x"0040";
    tmp(73753) := x"0040";
    tmp(73754) := x"0040";
    tmp(73755) := x"0040";
    tmp(73756) := x"0040";
    tmp(73757) := x"0840";
    tmp(73758) := x"0840";
    tmp(73759) := x"0840";
    tmp(73760) := x"0820";
    tmp(73761) := x"1020";
    tmp(73762) := x"1000";
    tmp(73763) := x"1800";
    tmp(73764) := x"1800";
    tmp(73765) := x"2020";
    tmp(73766) := x"2000";
    tmp(73767) := x"2000";
    tmp(73768) := x"2020";
    tmp(73769) := x"2020";
    tmp(73770) := x"2820";
    tmp(73771) := x"2820";
    tmp(73772) := x"2820";
    tmp(73773) := x"2000";
    tmp(73774) := x"2000";
    tmp(73775) := x"1800";
    tmp(73776) := x"2000";
    tmp(73777) := x"2820";
    tmp(73778) := x"3020";
    tmp(73779) := x"3020";
    tmp(73780) := x"3020";
    tmp(73781) := x"3820";
    tmp(73782) := x"3820";
    tmp(73783) := x"3020";
    tmp(73784) := x"3020";
    tmp(73785) := x"3020";
    tmp(73786) := x"3020";
    tmp(73787) := x"3820";
    tmp(73788) := x"2820";
    tmp(73789) := x"1800";
    tmp(73790) := x"1000";
    tmp(73791) := x"1800";
    tmp(73792) := x"2800";
    tmp(73793) := x"2800";
    tmp(73794) := x"2800";
    tmp(73795) := x"2000";
    tmp(73796) := x"1820";
    tmp(73797) := x"0820";
    tmp(73798) := x"0020";
    tmp(73799) := x"0020";
    tmp(73800) := x"0020";
    tmp(73801) := x"0020";
    tmp(73802) := x"0020";
    tmp(73803) := x"0820";
    tmp(73804) := x"0820";
    tmp(73805) := x"0820";
    tmp(73806) := x"0820";
    tmp(73807) := x"0820";
    tmp(73808) := x"0840";
    tmp(73809) := x"0840";
    tmp(73810) := x"0840";
    tmp(73811) := x"0840";
    tmp(73812) := x"0840";
    tmp(73813) := x"0840";
    tmp(73814) := x"0840";
    tmp(73815) := x"0840";
    tmp(73816) := x"0841";
    tmp(73817) := x"0840";
    tmp(73818) := x"0840";
    tmp(73819) := x"0841";
    tmp(73820) := x"0841";
    tmp(73821) := x"0840";
    tmp(73822) := x"0840";
    tmp(73823) := x"0840";
    tmp(73824) := x"0840";
    tmp(73825) := x"0840";
    tmp(73826) := x"0840";
    tmp(73827) := x"0840";
    tmp(73828) := x"0840";
    tmp(73829) := x"0840";
    tmp(73830) := x"0840";
    tmp(73831) := x"0840";
    tmp(73832) := x"0840";
    tmp(73833) := x"0840";
    tmp(73834) := x"0840";
    tmp(73835) := x"0840";
    tmp(73836) := x"0820";
    tmp(73837) := x"0820";
    tmp(73838) := x"0820";
    tmp(73839) := x"0820";
    tmp(73840) := x"0820";
    tmp(73841) := x"0820";
    tmp(73842) := x"0820";
    tmp(73843) := x"0820";
    tmp(73844) := x"0020";
    tmp(73845) := x"0020";
    tmp(73846) := x"0020";
    tmp(73847) := x"0020";
    tmp(73848) := x"0020";
    tmp(73849) := x"0020";
    tmp(73850) := x"0000";
    tmp(73851) := x"0020";
    tmp(73852) := x"0000";
    tmp(73853) := x"0000";
    tmp(73854) := x"0000";
    tmp(73855) := x"0000";
    tmp(73856) := x"0000";
    tmp(73857) := x"0000";
    tmp(73858) := x"0000";
    tmp(73859) := x"0000";
    tmp(73860) := x"0000";
    tmp(73861) := x"0000";
    tmp(73862) := x"0000";
    tmp(73863) := x"0000";
    tmp(73864) := x"0000";
    tmp(73865) := x"0020";
    tmp(73866) := x"0000";
    tmp(73867) := x"0000";
    tmp(73868) := x"0000";
    tmp(73869) := x"0000";
    tmp(73870) := x"0000";
    tmp(73871) := x"0000";
    tmp(73872) := x"0000";
    tmp(73873) := x"0000";
    tmp(73874) := x"0000";
    tmp(73875) := x"0000";
    tmp(73876) := x"0000";
    tmp(73877) := x"0000";
    tmp(73878) := x"0000";
    tmp(73879) := x"0000";
    tmp(73880) := x"0000";
    tmp(73881) := x"0020";
    tmp(73882) := x"0020";
    tmp(73883) := x"0020";
    tmp(73884) := x"0020";
    tmp(73885) := x"0020";
    tmp(73886) := x"0020";
    tmp(73887) := x"0020";
    tmp(73888) := x"0020";
    tmp(73889) := x"0020";
    tmp(73890) := x"0020";
    tmp(73891) := x"0020";
    tmp(73892) := x"0020";
    tmp(73893) := x"0020";
    tmp(73894) := x"0020";
    tmp(73895) := x"0020";
    tmp(73896) := x"0020";
    tmp(73897) := x"0020";
    tmp(73898) := x"0000";
    tmp(73899) := x"0020";
    tmp(73900) := x"0000";
    tmp(73901) := x"0000";
    tmp(73902) := x"0000";
    tmp(73903) := x"0000";
    tmp(73904) := x"0000";
    tmp(73905) := x"0000";
    tmp(73906) := x"0000";
    tmp(73907) := x"0000";
    tmp(73908) := x"0000";
    tmp(73909) := x"0000";
    tmp(73910) := x"0000";
    tmp(73911) := x"0000";
    tmp(73912) := x"0000";
    tmp(73913) := x"0000";
    tmp(73914) := x"0000";
    tmp(73915) := x"0000";
    tmp(73916) := x"0000";
    tmp(73917) := x"0000";
    tmp(73918) := x"0020";
    tmp(73919) := x"0000";
    tmp(73920) := x"0000";
    tmp(73921) := x"0020";
    tmp(73922) := x"0020";
    tmp(73923) := x"0020";
    tmp(73924) := x"0000";
    tmp(73925) := x"0020";
    tmp(73926) := x"0020";
    tmp(73927) := x"0020";
    tmp(73928) := x"0020";
    tmp(73929) := x"0020";
    tmp(73930) := x"0020";
    tmp(73931) := x"0020";
    tmp(73932) := x"0020";
    tmp(73933) := x"0020";
    tmp(73934) := x"0020";
    tmp(73935) := x"0020";
    tmp(73936) := x"0021";
    tmp(73937) := x"0021";
    tmp(73938) := x"0021";
    tmp(73939) := x"0041";
    tmp(73940) := x"0041";
    tmp(73941) := x"0041";
    tmp(73942) := x"0061";
    tmp(73943) := x"0081";
    tmp(73944) := x"0081";
    tmp(73945) := x"0081";
    tmp(73946) := x"0061";
    tmp(73947) := x"0061";
    tmp(73948) := x"0061";
    tmp(73949) := x"0061";
    tmp(73950) := x"0061";
    tmp(73951) := x"0061";
    tmp(73952) := x"0061";
    tmp(73953) := x"0061";
    tmp(73954) := x"0060";
    tmp(73955) := x"0040";
    tmp(73956) := x"0040";
    tmp(73957) := x"0040";
    tmp(73958) := x"0020";
    tmp(73959) := x"0040";
    tmp(73960) := x"0041";
    tmp(73961) := x"0041";
    tmp(73962) := x"0041";
    tmp(73963) := x"0040";
    tmp(73964) := x"0040";
    tmp(73965) := x"0040";
    tmp(73966) := x"0040";
    tmp(73967) := x"0040";
    tmp(73968) := x"0040";
    tmp(73969) := x"0040";
    tmp(73970) := x"0040";
    tmp(73971) := x"0040";
    tmp(73972) := x"0020";
    tmp(73973) := x"0020";
    tmp(73974) := x"0020";
    tmp(73975) := x"0020";
    tmp(73976) := x"0040";
    tmp(73977) := x"0040";
    tmp(73978) := x"0060";
    tmp(73979) := x"0860";
    tmp(73980) := x"0040";
    tmp(73981) := x"0020";
    tmp(73982) := x"0020";
    tmp(73983) := x"0020";
    tmp(73984) := x"0020";
    tmp(73985) := x"0020";
    tmp(73986) := x"0020";
    tmp(73987) := x"0020";
    tmp(73988) := x"0040";
    tmp(73989) := x"0040";
    tmp(73990) := x"0040";
    tmp(73991) := x"0040";
    tmp(73992) := x"0040";
    tmp(73993) := x"0040";
    tmp(73994) := x"0840";
    tmp(73995) := x"0820";
    tmp(73996) := x"0820";
    tmp(73997) := x"0820";
    tmp(73998) := x"0820";
    tmp(73999) := x"0820";
    tmp(74000) := x"1020";
    tmp(74001) := x"1000";
    tmp(74002) := x"1000";
    tmp(74003) := x"1800";
    tmp(74004) := x"2000";
    tmp(74005) := x"2820";
    tmp(74006) := x"2820";
    tmp(74007) := x"2820";
    tmp(74008) := x"2820";
    tmp(74009) := x"1800";
    tmp(74010) := x"2000";
    tmp(74011) := x"2820";
    tmp(74012) := x"2800";
    tmp(74013) := x"3000";
    tmp(74014) := x"3020";
    tmp(74015) := x"2800";
    tmp(74016) := x"3020";
    tmp(74017) := x"3820";
    tmp(74018) := x"3820";
    tmp(74019) := x"3820";
    tmp(74020) := x"3820";
    tmp(74021) := x"3020";
    tmp(74022) := x"3020";
    tmp(74023) := x"3020";
    tmp(74024) := x"3020";
    tmp(74025) := x"3020";
    tmp(74026) := x"2820";
    tmp(74027) := x"2000";
    tmp(74028) := x"1000";
    tmp(74029) := x"0800";
    tmp(74030) := x"1800";
    tmp(74031) := x"2800";
    tmp(74032) := x"2800";
    tmp(74033) := x"2800";
    tmp(74034) := x"2000";
    tmp(74035) := x"1800";
    tmp(74036) := x"0820";
    tmp(74037) := x"0820";
    tmp(74038) := x"0020";
    tmp(74039) := x"0020";
    tmp(74040) := x"0020";
    tmp(74041) := x"0020";
    tmp(74042) := x"0020";
    tmp(74043) := x"0020";
    tmp(74044) := x"0020";
    tmp(74045) := x"0020";
    tmp(74046) := x"0820";
    tmp(74047) := x"0820";
    tmp(74048) := x"0820";
    tmp(74049) := x"0820";
    tmp(74050) := x"0820";
    tmp(74051) := x"0820";
    tmp(74052) := x"0840";
    tmp(74053) := x"0840";
    tmp(74054) := x"0840";
    tmp(74055) := x"0840";
    tmp(74056) := x"0840";
    tmp(74057) := x"0840";
    tmp(74058) := x"0840";
    tmp(74059) := x"0840";
    tmp(74060) := x"0840";
    tmp(74061) := x"0840";
    tmp(74062) := x"0840";
    tmp(74063) := x"0840";
    tmp(74064) := x"0840";
    tmp(74065) := x"0840";
    tmp(74066) := x"0840";
    tmp(74067) := x"0840";
    tmp(74068) := x"0840";
    tmp(74069) := x"0840";
    tmp(74070) := x"0840";
    tmp(74071) := x"0820";
    tmp(74072) := x"0820";
    tmp(74073) := x"0820";
    tmp(74074) := x"0820";
    tmp(74075) := x"0820";
    tmp(74076) := x"0820";
    tmp(74077) := x"0820";
    tmp(74078) := x"0820";
    tmp(74079) := x"0820";
    tmp(74080) := x"0820";
    tmp(74081) := x"0020";
    tmp(74082) := x"0020";
    tmp(74083) := x"0020";
    tmp(74084) := x"0020";
    tmp(74085) := x"0020";
    tmp(74086) := x"0020";
    tmp(74087) := x"0000";
    tmp(74088) := x"0020";
    tmp(74089) := x"0000";
    tmp(74090) := x"0000";
    tmp(74091) := x"0000";
    tmp(74092) := x"0000";
    tmp(74093) := x"0000";
    tmp(74094) := x"0000";
    tmp(74095) := x"0000";
    tmp(74096) := x"0000";
    tmp(74097) := x"0000";
    tmp(74098) := x"0000";
    tmp(74099) := x"0000";
    tmp(74100) := x"0000";
    tmp(74101) := x"0000";
    tmp(74102) := x"0000";
    tmp(74103) := x"0000";
    tmp(74104) := x"0000";
    tmp(74105) := x"0000";
    tmp(74106) := x"0000";
    tmp(74107) := x"0000";
    tmp(74108) := x"0000";
    tmp(74109) := x"0000";
    tmp(74110) := x"0020";
    tmp(74111) := x"0000";
    tmp(74112) := x"0000";
    tmp(74113) := x"0000";
    tmp(74114) := x"0000";
    tmp(74115) := x"0000";
    tmp(74116) := x"0000";
    tmp(74117) := x"0000";
    tmp(74118) := x"0000";
    tmp(74119) := x"0000";
    tmp(74120) := x"0000";
    tmp(74121) := x"0000";
    tmp(74122) := x"0000";
    tmp(74123) := x"0000";
    tmp(74124) := x"0000";
    tmp(74125) := x"0000";
    tmp(74126) := x"0020";
    tmp(74127) := x"0020";
    tmp(74128) := x"0020";
    tmp(74129) := x"0020";
    tmp(74130) := x"0020";
    tmp(74131) := x"0020";
    tmp(74132) := x"0020";
    tmp(74133) := x"0020";
    tmp(74134) := x"0000";
    tmp(74135) := x"0000";
    tmp(74136) := x"0000";
    tmp(74137) := x"0000";
    tmp(74138) := x"0000";
    tmp(74139) := x"0000";
    tmp(74140) := x"0000";
    tmp(74141) := x"0000";
    tmp(74142) := x"0000";
    tmp(74143) := x"0000";
    tmp(74144) := x"0000";
    tmp(74145) := x"0000";
    tmp(74146) := x"0000";
    tmp(74147) := x"0000";
    tmp(74148) := x"0000";
    tmp(74149) := x"0000";
    tmp(74150) := x"0000";
    tmp(74151) := x"0000";
    tmp(74152) := x"0000";
    tmp(74153) := x"0000";
    tmp(74154) := x"0000";
    tmp(74155) := x"0000";
    tmp(74156) := x"0000";
    tmp(74157) := x"0000";
    tmp(74158) := x"0000";
    tmp(74159) := x"0020";
    tmp(74160) := x"0000";
    tmp(74161) := x"0020";
    tmp(74162) := x"0020";
    tmp(74163) := x"0020";
    tmp(74164) := x"0020";
    tmp(74165) := x"0020";
    tmp(74166) := x"0020";
    tmp(74167) := x"0021";
    tmp(74168) := x"0021";
    tmp(74169) := x"0021";
    tmp(74170) := x"0021";
    tmp(74171) := x"0020";
    tmp(74172) := x"0020";
    tmp(74173) := x"0020";
    tmp(74174) := x"0020";
    tmp(74175) := x"0020";
    tmp(74176) := x"0020";
    tmp(74177) := x"0020";
    tmp(74178) := x"0020";
    tmp(74179) := x"0020";
    tmp(74180) := x"0020";
    tmp(74181) := x"0020";
    tmp(74182) := x"0020";
    tmp(74183) := x"0020";
    tmp(74184) := x"0041";
    tmp(74185) := x"0041";
    tmp(74186) := x"0061";
    tmp(74187) := x"0061";
    tmp(74188) := x"0081";
    tmp(74189) := x"0081";
    tmp(74190) := x"0081";
    tmp(74191) := x"0061";
    tmp(74192) := x"0061";
    tmp(74193) := x"0041";
    tmp(74194) := x"0060";
    tmp(74195) := x"0060";
    tmp(74196) := x"0040";
    tmp(74197) := x"0040";
    tmp(74198) := x"0040";
    tmp(74199) := x"0040";
    tmp(74200) := x"0041";
    tmp(74201) := x"0081";
    tmp(74202) := x"0061";
    tmp(74203) := x"0061";
    tmp(74204) := x"0041";
    tmp(74205) := x"0040";
    tmp(74206) := x"0040";
    tmp(74207) := x"0040";
    tmp(74208) := x"0040";
    tmp(74209) := x"0040";
    tmp(74210) := x"0040";
    tmp(74211) := x"0040";
    tmp(74212) := x"0041";
    tmp(74213) := x"0041";
    tmp(74214) := x"0040";
    tmp(74215) := x"0040";
    tmp(74216) := x"0040";
    tmp(74217) := x"0040";
    tmp(74218) := x"0840";
    tmp(74219) := x"0040";
    tmp(74220) := x"0040";
    tmp(74221) := x"0020";
    tmp(74222) := x"0020";
    tmp(74223) := x"0000";
    tmp(74224) := x"0020";
    tmp(74225) := x"0020";
    tmp(74226) := x"0020";
    tmp(74227) := x"0020";
    tmp(74228) := x"0040";
    tmp(74229) := x"0840";
    tmp(74230) := x"0840";
    tmp(74231) := x"0840";
    tmp(74232) := x"0840";
    tmp(74233) := x"0820";
    tmp(74234) := x"0820";
    tmp(74235) := x"0800";
    tmp(74236) := x"0800";
    tmp(74237) := x"1000";
    tmp(74238) := x"1000";
    tmp(74239) := x"1000";
    tmp(74240) := x"1000";
    tmp(74241) := x"1000";
    tmp(74242) := x"1000";
    tmp(74243) := x"1800";
    tmp(74244) := x"1800";
    tmp(74245) := x"2800";
    tmp(74246) := x"2820";
    tmp(74247) := x"2800";
    tmp(74248) := x"1800";
    tmp(74249) := x"1000";
    tmp(74250) := x"2020";
    tmp(74251) := x"2820";
    tmp(74252) := x"3020";
    tmp(74253) := x"3820";
    tmp(74254) := x"3020";
    tmp(74255) := x"3020";
    tmp(74256) := x"3020";
    tmp(74257) := x"3020";
    tmp(74258) := x"3020";
    tmp(74259) := x"2820";
    tmp(74260) := x"2800";
    tmp(74261) := x"2000";
    tmp(74262) := x"2800";
    tmp(74263) := x"2800";
    tmp(74264) := x"2800";
    tmp(74265) := x"2800";
    tmp(74266) := x"1800";
    tmp(74267) := x"1000";
    tmp(74268) := x"0800";
    tmp(74269) := x"0800";
    tmp(74270) := x"3020";
    tmp(74271) := x"2800";
    tmp(74272) := x"2000";
    tmp(74273) := x"2000";
    tmp(74274) := x"1800";
    tmp(74275) := x"1020";
    tmp(74276) := x"0820";
    tmp(74277) := x"0020";
    tmp(74278) := x"0020";
    tmp(74279) := x"0020";
    tmp(74280) := x"0020";
    tmp(74281) := x"0020";
    tmp(74282) := x"0020";
    tmp(74283) := x"0020";
    tmp(74284) := x"0020";
    tmp(74285) := x"0020";
    tmp(74286) := x"0020";
    tmp(74287) := x"0020";
    tmp(74288) := x"0820";
    tmp(74289) := x"0820";
    tmp(74290) := x"0820";
    tmp(74291) := x"0820";
    tmp(74292) := x"0820";
    tmp(74293) := x"0820";
    tmp(74294) := x"0820";
    tmp(74295) := x"0820";
    tmp(74296) := x"0820";
    tmp(74297) := x"0840";
    tmp(74298) := x"0840";
    tmp(74299) := x"0840";
    tmp(74300) := x"0840";
    tmp(74301) := x"0840";
    tmp(74302) := x"0840";
    tmp(74303) := x"0840";
    tmp(74304) := x"0840";
    tmp(74305) := x"0840";
    tmp(74306) := x"0840";
    tmp(74307) := x"0820";
    tmp(74308) := x"0820";
    tmp(74309) := x"0820";
    tmp(74310) := x"0820";
    tmp(74311) := x"0820";
    tmp(74312) := x"0820";
    tmp(74313) := x"0820";
    tmp(74314) := x"0820";
    tmp(74315) := x"0820";
    tmp(74316) := x"0820";
    tmp(74317) := x"0820";
    tmp(74318) := x"0820";
    tmp(74319) := x"0020";
    tmp(74320) := x"0020";
    tmp(74321) := x"0020";
    tmp(74322) := x"0020";
    tmp(74323) := x"0020";
    tmp(74324) := x"0020";
    tmp(74325) := x"0020";
    tmp(74326) := x"0000";
    tmp(74327) := x"0020";
    tmp(74328) := x"0000";
    tmp(74329) := x"0000";
    tmp(74330) := x"0000";
    tmp(74331) := x"0000";
    tmp(74332) := x"0020";
    tmp(74333) := x"0000";
    tmp(74334) := x"0000";
    tmp(74335) := x"0000";
    tmp(74336) := x"0000";
    tmp(74337) := x"0000";
    tmp(74338) := x"0000";
    tmp(74339) := x"0000";
    tmp(74340) := x"0000";
    tmp(74341) := x"0000";
    tmp(74342) := x"0000";
    tmp(74343) := x"0000";
    tmp(74344) := x"0000";
    tmp(74345) := x"0000";
    tmp(74346) := x"0000";
    tmp(74347) := x"0000";
    tmp(74348) := x"0000";
    tmp(74349) := x"0000";
    tmp(74350) := x"0000";
    tmp(74351) := x"0000";
    tmp(74352) := x"0000";
    tmp(74353) := x"0000";
    tmp(74354) := x"0000";
    tmp(74355) := x"0000";
    tmp(74356) := x"0000";
    tmp(74357) := x"0000";
    tmp(74358) := x"0000";
    tmp(74359) := x"0000";
    tmp(74360) := x"0000";
    tmp(74361) := x"0000";
    tmp(74362) := x"0000";
    tmp(74363) := x"0000";
    tmp(74364) := x"0000";
    tmp(74365) := x"0000";
    tmp(74366) := x"0000";
    tmp(74367) := x"0000";
    tmp(74368) := x"0000";
    tmp(74369) := x"0000";
    tmp(74370) := x"0000";
    tmp(74371) := x"0000";
    tmp(74372) := x"0000";
    tmp(74373) := x"0000";
    tmp(74374) := x"0000";
    tmp(74375) := x"0000";
    tmp(74376) := x"0000";
    tmp(74377) := x"0000";
    tmp(74378) := x"0000";
    tmp(74379) := x"0000";
    tmp(74380) := x"0000";
    tmp(74381) := x"0000";
    tmp(74382) := x"0000";
    tmp(74383) := x"0000";
    tmp(74384) := x"0000";
    tmp(74385) := x"0000";
    tmp(74386) := x"0000";
    tmp(74387) := x"0000";
    tmp(74388) := x"0000";
    tmp(74389) := x"0000";
    tmp(74390) := x"0000";
    tmp(74391) := x"0000";
    tmp(74392) := x"0000";
    tmp(74393) := x"0000";
    tmp(74394) := x"0000";
    tmp(74395) := x"0000";
    tmp(74396) := x"0000";
    tmp(74397) := x"0000";
    tmp(74398) := x"0020";
    tmp(74399) := x"0020";
    tmp(74400) := x"0000";
    tmp(74401) := x"0000";
    tmp(74402) := x"0000";
    tmp(74403) := x"0000";
    tmp(74404) := x"0020";
    tmp(74405) := x"0000";
    tmp(74406) := x"0020";
    tmp(74407) := x"0020";
    tmp(74408) := x"0021";
    tmp(74409) := x"0041";
    tmp(74410) := x"0041";
    tmp(74411) := x"0041";
    tmp(74412) := x"0020";
    tmp(74413) := x"0020";
    tmp(74414) := x"0020";
    tmp(74415) := x"0020";
    tmp(74416) := x"0020";
    tmp(74417) := x"0020";
    tmp(74418) := x"0020";
    tmp(74419) := x"0020";
    tmp(74420) := x"0020";
    tmp(74421) := x"0020";
    tmp(74422) := x"0020";
    tmp(74423) := x"0020";
    tmp(74424) := x"0020";
    tmp(74425) := x"0020";
    tmp(74426) := x"0020";
    tmp(74427) := x"0020";
    tmp(74428) := x"0020";
    tmp(74429) := x"0041";
    tmp(74430) := x"0041";
    tmp(74431) := x"0041";
    tmp(74432) := x"0040";
    tmp(74433) := x"0040";
    tmp(74434) := x"0040";
    tmp(74435) := x"0040";
    tmp(74436) := x"0060";
    tmp(74437) := x"0040";
    tmp(74438) := x"0040";
    tmp(74439) := x"0040";
    tmp(74440) := x"0040";
    tmp(74441) := x"0040";
    tmp(74442) := x"0061";
    tmp(74443) := x"0881";
    tmp(74444) := x"0061";
    tmp(74445) := x"0061";
    tmp(74446) := x"0041";
    tmp(74447) := x"0041";
    tmp(74448) := x"0040";
    tmp(74449) := x"0040";
    tmp(74450) := x"0040";
    tmp(74451) := x"0040";
    tmp(74452) := x"0041";
    tmp(74453) := x"0020";
    tmp(74454) := x"0040";
    tmp(74455) := x"0040";
    tmp(74456) := x"0040";
    tmp(74457) := x"0040";
    tmp(74458) := x"0040";
    tmp(74459) := x"0020";
    tmp(74460) := x"0040";
    tmp(74461) := x"0020";
    tmp(74462) := x"0020";
    tmp(74463) := x"0020";
    tmp(74464) := x"0020";
    tmp(74465) := x"0020";
    tmp(74466) := x"0020";
    tmp(74467) := x"0020";
    tmp(74468) := x"0020";
    tmp(74469) := x"0020";
    tmp(74470) := x"0020";
    tmp(74471) := x"0820";
    tmp(74472) := x"0820";
    tmp(74473) := x"0800";
    tmp(74474) := x"0800";
    tmp(74475) := x"0800";
    tmp(74476) := x"0800";
    tmp(74477) := x"0800";
    tmp(74478) := x"0800";
    tmp(74479) := x"0800";
    tmp(74480) := x"0800";
    tmp(74481) := x"0800";
    tmp(74482) := x"0800";
    tmp(74483) := x"1000";
    tmp(74484) := x"2000";
    tmp(74485) := x"2000";
    tmp(74486) := x"2000";
    tmp(74487) := x"2000";
    tmp(74488) := x"1800";
    tmp(74489) := x"1820";
    tmp(74490) := x"2020";
    tmp(74491) := x"2820";
    tmp(74492) := x"3820";
    tmp(74493) := x"3020";
    tmp(74494) := x"3000";
    tmp(74495) := x"3020";
    tmp(74496) := x"3020";
    tmp(74497) := x"2000";
    tmp(74498) := x"2000";
    tmp(74499) := x"2820";
    tmp(74500) := x"2820";
    tmp(74501) := x"2820";
    tmp(74502) := x"2800";
    tmp(74503) := x"3020";
    tmp(74504) := x"3020";
    tmp(74505) := x"2800";
    tmp(74506) := x"2000";
    tmp(74507) := x"1800";
    tmp(74508) := x"1000";
    tmp(74509) := x"1000";
    tmp(74510) := x"3020";
    tmp(74511) := x"1800";
    tmp(74512) := x"1800";
    tmp(74513) := x"1800";
    tmp(74514) := x"1820";
    tmp(74515) := x"0820";
    tmp(74516) := x"0020";
    tmp(74517) := x"0020";
    tmp(74518) := x"0020";
    tmp(74519) := x"0020";
    tmp(74520) := x"0020";
    tmp(74521) := x"0020";
    tmp(74522) := x"0020";
    tmp(74523) := x"0020";
    tmp(74524) := x"0020";
    tmp(74525) := x"0020";
    tmp(74526) := x"0020";
    tmp(74527) := x"0020";
    tmp(74528) := x"0020";
    tmp(74529) := x"0020";
    tmp(74530) := x"0020";
    tmp(74531) := x"0020";
    tmp(74532) := x"0020";
    tmp(74533) := x"0820";
    tmp(74534) := x"0820";
    tmp(74535) := x"0820";
    tmp(74536) := x"0820";
    tmp(74537) := x"0820";
    tmp(74538) := x"0820";
    tmp(74539) := x"0820";
    tmp(74540) := x"0820";
    tmp(74541) := x"0820";
    tmp(74542) := x"0820";
    tmp(74543) := x"0820";
    tmp(74544) := x"0820";
    tmp(74545) := x"0820";
    tmp(74546) := x"0820";
    tmp(74547) := x"0820";
    tmp(74548) := x"0820";
    tmp(74549) := x"0820";
    tmp(74550) := x"0820";
    tmp(74551) := x"0820";
    tmp(74552) := x"0820";
    tmp(74553) := x"0820";
    tmp(74554) := x"0820";
    tmp(74555) := x"0820";
    tmp(74556) := x"0820";
    tmp(74557) := x"0020";
    tmp(74558) := x"0020";
    tmp(74559) := x"0020";
    tmp(74560) := x"0020";
    tmp(74561) := x"0020";
    tmp(74562) := x"0020";
    tmp(74563) := x"0020";
    tmp(74564) := x"0020";
    tmp(74565) := x"0020";
    tmp(74566) := x"0020";
    tmp(74567) := x"0000";
    tmp(74568) := x"0000";
    tmp(74569) := x"0000";
    tmp(74570) := x"0000";
    tmp(74571) := x"0020";
    tmp(74572) := x"0000";
    tmp(74573) := x"0000";
    tmp(74574) := x"0000";
    tmp(74575) := x"0000";
    tmp(74576) := x"0000";
    tmp(74577) := x"0000";
    tmp(74578) := x"0000";
    tmp(74579) := x"0000";
    tmp(74580) := x"0000";
    tmp(74581) := x"0000";
    tmp(74582) := x"0000";
    tmp(74583) := x"0000";
    tmp(74584) := x"0000";
    tmp(74585) := x"0000";
    tmp(74586) := x"0000";
    tmp(74587) := x"0000";
    tmp(74588) := x"0000";
    tmp(74589) := x"0000";
    tmp(74590) := x"0000";
    tmp(74591) := x"0000";
    tmp(74592) := x"0000";
    tmp(74593) := x"0000";
    tmp(74594) := x"0000";
    tmp(74595) := x"0000";
    tmp(74596) := x"0000";
    tmp(74597) := x"0000";
    tmp(74598) := x"0000";
    tmp(74599) := x"0000";
    tmp(74600) := x"0000";
    tmp(74601) := x"0000";
    tmp(74602) := x"0000";
    tmp(74603) := x"0000";
    tmp(74604) := x"0000";
    tmp(74605) := x"0000";
    tmp(74606) := x"0000";
    tmp(74607) := x"0000";
    tmp(74608) := x"0000";
    tmp(74609) := x"0000";
    tmp(74610) := x"0000";
    tmp(74611) := x"0000";
    tmp(74612) := x"0000";
    tmp(74613) := x"0000";
    tmp(74614) := x"0000";
    tmp(74615) := x"0000";
    tmp(74616) := x"0000";
    tmp(74617) := x"0000";
    tmp(74618) := x"0000";
    tmp(74619) := x"0000";
    tmp(74620) := x"0000";
    tmp(74621) := x"0000";
    tmp(74622) := x"0000";
    tmp(74623) := x"0000";
    tmp(74624) := x"0000";
    tmp(74625) := x"0000";
    tmp(74626) := x"0000";
    tmp(74627) := x"0000";
    tmp(74628) := x"0000";
    tmp(74629) := x"0000";
    tmp(74630) := x"0000";
    tmp(74631) := x"0000";
    tmp(74632) := x"0000";
    tmp(74633) := x"0000";
    tmp(74634) := x"0000";
    tmp(74635) := x"0000";
    tmp(74636) := x"0000";
    tmp(74637) := x"0000";
    tmp(74638) := x"0020";
    tmp(74639) := x"0020";
    tmp(74640) := x"0000";
    tmp(74641) := x"0000";
    tmp(74642) := x"0000";
    tmp(74643) := x"0000";
    tmp(74644) := x"0000";
    tmp(74645) := x"0000";
    tmp(74646) := x"0000";
    tmp(74647) := x"0000";
    tmp(74648) := x"0020";
    tmp(74649) := x"0021";
    tmp(74650) := x"0041";
    tmp(74651) := x"0041";
    tmp(74652) := x"0021";
    tmp(74653) := x"0020";
    tmp(74654) := x"0020";
    tmp(74655) := x"0020";
    tmp(74656) := x"0020";
    tmp(74657) := x"0020";
    tmp(74658) := x"0020";
    tmp(74659) := x"0020";
    tmp(74660) := x"0020";
    tmp(74661) := x"0020";
    tmp(74662) := x"0020";
    tmp(74663) := x"0020";
    tmp(74664) := x"0020";
    tmp(74665) := x"0020";
    tmp(74666) := x"0020";
    tmp(74667) := x"0020";
    tmp(74668) := x"0020";
    tmp(74669) := x"0020";
    tmp(74670) := x"0020";
    tmp(74671) := x"0020";
    tmp(74672) := x"0040";
    tmp(74673) := x"0040";
    tmp(74674) := x"0040";
    tmp(74675) := x"0040";
    tmp(74676) := x"0040";
    tmp(74677) := x"0040";
    tmp(74678) := x"0060";
    tmp(74679) := x"0060";
    tmp(74680) := x"0040";
    tmp(74681) := x"0040";
    tmp(74682) := x"0041";
    tmp(74683) := x"0041";
    tmp(74684) := x"0061";
    tmp(74685) := x"0881";
    tmp(74686) := x"0881";
    tmp(74687) := x"0061";
    tmp(74688) := x"0060";
    tmp(74689) := x"0060";
    tmp(74690) := x"0040";
    tmp(74691) := x"0040";
    tmp(74692) := x"0040";
    tmp(74693) := x"0020";
    tmp(74694) := x"0020";
    tmp(74695) := x"0020";
    tmp(74696) := x"0040";
    tmp(74697) := x"0040";
    tmp(74698) := x"0020";
    tmp(74699) := x"0040";
    tmp(74700) := x"0040";
    tmp(74701) := x"0020";
    tmp(74702) := x"0020";
    tmp(74703) := x"0020";
    tmp(74704) := x"0020";
    tmp(74705) := x"0020";
    tmp(74706) := x"0020";
    tmp(74707) := x"0020";
    tmp(74708) := x"0020";
    tmp(74709) := x"0020";
    tmp(74710) := x"0820";
    tmp(74711) := x"0820";
    tmp(74712) := x"0820";
    tmp(74713) := x"0800";
    tmp(74714) := x"0800";
    tmp(74715) := x"0800";
    tmp(74716) := x"0800";
    tmp(74717) := x"0800";
    tmp(74718) := x"1000";
    tmp(74719) := x"1000";
    tmp(74720) := x"1000";
    tmp(74721) := x"1000";
    tmp(74722) := x"1000";
    tmp(74723) := x"1800";
    tmp(74724) := x"2000";
    tmp(74725) := x"2000";
    tmp(74726) := x"2000";
    tmp(74727) := x"2000";
    tmp(74728) := x"2000";
    tmp(74729) := x"2000";
    tmp(74730) := x"2800";
    tmp(74731) := x"2820";
    tmp(74732) := x"2820";
    tmp(74733) := x"2800";
    tmp(74734) := x"3000";
    tmp(74735) := x"3020";
    tmp(74736) := x"2800";
    tmp(74737) := x"2000";
    tmp(74738) := x"2800";
    tmp(74739) := x"2820";
    tmp(74740) := x"2820";
    tmp(74741) := x"2800";
    tmp(74742) := x"2820";
    tmp(74743) := x"2820";
    tmp(74744) := x"3020";
    tmp(74745) := x"3020";
    tmp(74746) := x"2820";
    tmp(74747) := x"1800";
    tmp(74748) := x"0800";
    tmp(74749) := x"2000";
    tmp(74750) := x"2000";
    tmp(74751) := x"1000";
    tmp(74752) := x"1820";
    tmp(74753) := x"1820";
    tmp(74754) := x"0820";
    tmp(74755) := x"0020";
    tmp(74756) := x"0020";
    tmp(74757) := x"0000";
    tmp(74758) := x"0000";
    tmp(74759) := x"0000";
    tmp(74760) := x"0000";
    tmp(74761) := x"0000";
    tmp(74762) := x"0000";
    tmp(74763) := x"0020";
    tmp(74764) := x"0000";
    tmp(74765) := x"0020";
    tmp(74766) := x"0020";
    tmp(74767) := x"0020";
    tmp(74768) := x"0020";
    tmp(74769) := x"0020";
    tmp(74770) := x"0020";
    tmp(74771) := x"0020";
    tmp(74772) := x"0020";
    tmp(74773) := x"0020";
    tmp(74774) := x"0020";
    tmp(74775) := x"0820";
    tmp(74776) := x"0820";
    tmp(74777) := x"0820";
    tmp(74778) := x"0820";
    tmp(74779) := x"0820";
    tmp(74780) := x"0820";
    tmp(74781) := x"0820";
    tmp(74782) := x"0820";
    tmp(74783) := x"0820";
    tmp(74784) := x"0820";
    tmp(74785) := x"0820";
    tmp(74786) := x"0820";
    tmp(74787) := x"0820";
    tmp(74788) := x"0820";
    tmp(74789) := x"0820";
    tmp(74790) := x"0820";
    tmp(74791) := x"0820";
    tmp(74792) := x"0020";
    tmp(74793) := x"0020";
    tmp(74794) := x"0020";
    tmp(74795) := x"0020";
    tmp(74796) := x"0020";
    tmp(74797) := x"0020";
    tmp(74798) := x"0020";
    tmp(74799) := x"0020";
    tmp(74800) := x"0020";
    tmp(74801) := x"0020";
    tmp(74802) := x"0020";
    tmp(74803) := x"0020";
    tmp(74804) := x"0020";
    tmp(74805) := x"0000";
    tmp(74806) := x"0020";
    tmp(74807) := x"0020";
    tmp(74808) := x"0000";
    tmp(74809) := x"0000";
    tmp(74810) := x"0000";
    tmp(74811) := x"0000";
    tmp(74812) := x"0000";
    tmp(74813) := x"0000";
    tmp(74814) := x"0000";
    tmp(74815) := x"0000";
    tmp(74816) := x"0000";
    tmp(74817) := x"0000";
    tmp(74818) := x"0000";
    tmp(74819) := x"0000";
    tmp(74820) := x"0000";
    tmp(74821) := x"0000";
    tmp(74822) := x"0000";
    tmp(74823) := x"0000";
    tmp(74824) := x"0000";
    tmp(74825) := x"0000";
    tmp(74826) := x"0000";
    tmp(74827) := x"0000";
    tmp(74828) := x"0000";
    tmp(74829) := x"0000";
    tmp(74830) := x"0000";
    tmp(74831) := x"0000";
    tmp(74832) := x"0000";
    tmp(74833) := x"0000";
    tmp(74834) := x"0000";
    tmp(74835) := x"0000";
    tmp(74836) := x"0000";
    tmp(74837) := x"0000";
    tmp(74838) := x"0000";
    tmp(74839) := x"0000";
    tmp(74840) := x"0000";
    tmp(74841) := x"0000";
    tmp(74842) := x"0000";
    tmp(74843) := x"0000";
    tmp(74844) := x"0000";
    tmp(74845) := x"0000";
    tmp(74846) := x"0000";
    tmp(74847) := x"0000";
    tmp(74848) := x"0000";
    tmp(74849) := x"0000";
    tmp(74850) := x"0000";
    tmp(74851) := x"0000";
    tmp(74852) := x"0000";
    tmp(74853) := x"0000";
    tmp(74854) := x"0000";
    tmp(74855) := x"0000";
    tmp(74856) := x"0000";
    tmp(74857) := x"0000";
    tmp(74858) := x"0000";
    tmp(74859) := x"0000";
    tmp(74860) := x"0000";
    tmp(74861) := x"0000";
    tmp(74862) := x"0000";
    tmp(74863) := x"0000";
    tmp(74864) := x"0000";
    tmp(74865) := x"0000";
    tmp(74866) := x"0000";
    tmp(74867) := x"0000";
    tmp(74868) := x"0000";
    tmp(74869) := x"0000";
    tmp(74870) := x"0000";
    tmp(74871) := x"0000";
    tmp(74872) := x"0000";
    tmp(74873) := x"0000";
    tmp(74874) := x"0000";
    tmp(74875) := x"0000";
    tmp(74876) := x"0000";
    tmp(74877) := x"0000";
    tmp(74878) := x"0000";
    tmp(74879) := x"0000";
    tmp(74880) := x"0000";
    tmp(74881) := x"0000";
    tmp(74882) := x"0000";
    tmp(74883) := x"0000";
    tmp(74884) := x"0000";
    tmp(74885) := x"0000";
    tmp(74886) := x"0000";
    tmp(74887) := x"0000";
    tmp(74888) := x"0000";
    tmp(74889) := x"0000";
    tmp(74890) := x"0020";
    tmp(74891) := x"0041";
    tmp(74892) := x"0041";
    tmp(74893) := x"0041";
    tmp(74894) := x"0021";
    tmp(74895) := x"0020";
    tmp(74896) := x"0020";
    tmp(74897) := x"0020";
    tmp(74898) := x"0020";
    tmp(74899) := x"0020";
    tmp(74900) := x"0020";
    tmp(74901) := x"0020";
    tmp(74902) := x"0020";
    tmp(74903) := x"0020";
    tmp(74904) := x"0020";
    tmp(74905) := x"0020";
    tmp(74906) := x"0020";
    tmp(74907) := x"0020";
    tmp(74908) := x"0020";
    tmp(74909) := x"0020";
    tmp(74910) := x"0020";
    tmp(74911) := x"0040";
    tmp(74912) := x"0040";
    tmp(74913) := x"0040";
    tmp(74914) := x"0040";
    tmp(74915) := x"0040";
    tmp(74916) := x"0040";
    tmp(74917) := x"0040";
    tmp(74918) := x"0040";
    tmp(74919) := x"0040";
    tmp(74920) := x"0860";
    tmp(74921) := x"0060";
    tmp(74922) := x"0040";
    tmp(74923) := x"0041";
    tmp(74924) := x"0040";
    tmp(74925) := x"0040";
    tmp(74926) := x"0060";
    tmp(74927) := x"0060";
    tmp(74928) := x"0860";
    tmp(74929) := x"0060";
    tmp(74930) := x"0040";
    tmp(74931) := x"0040";
    tmp(74932) := x"0040";
    tmp(74933) := x"0020";
    tmp(74934) := x"0020";
    tmp(74935) := x"0020";
    tmp(74936) := x"0020";
    tmp(74937) := x"0020";
    tmp(74938) := x"0020";
    tmp(74939) := x"0040";
    tmp(74940) := x"0040";
    tmp(74941) := x"0020";
    tmp(74942) := x"0020";
    tmp(74943) := x"0020";
    tmp(74944) := x"0000";
    tmp(74945) := x"0000";
    tmp(74946) := x"0000";
    tmp(74947) := x"0000";
    tmp(74948) := x"0000";
    tmp(74949) := x"0020";
    tmp(74950) := x"0820";
    tmp(74951) := x"0820";
    tmp(74952) := x"0820";
    tmp(74953) := x"0800";
    tmp(74954) := x"0800";
    tmp(74955) := x"1000";
    tmp(74956) := x"1000";
    tmp(74957) := x"1800";
    tmp(74958) := x"1800";
    tmp(74959) := x"2000";
    tmp(74960) := x"1800";
    tmp(74961) := x"1800";
    tmp(74962) := x"1800";
    tmp(74963) := x"1800";
    tmp(74964) := x"2000";
    tmp(74965) := x"2820";
    tmp(74966) := x"2820";
    tmp(74967) := x"2820";
    tmp(74968) := x"2800";
    tmp(74969) := x"2800";
    tmp(74970) := x"2800";
    tmp(74971) := x"2820";
    tmp(74972) := x"2820";
    tmp(74973) := x"2800";
    tmp(74974) := x"2800";
    tmp(74975) := x"2800";
    tmp(74976) := x"2800";
    tmp(74977) := x"2800";
    tmp(74978) := x"2820";
    tmp(74979) := x"2820";
    tmp(74980) := x"2820";
    tmp(74981) := x"2820";
    tmp(74982) := x"2020";
    tmp(74983) := x"2020";
    tmp(74984) := x"1800";
    tmp(74985) := x"1800";
    tmp(74986) := x"0800";
    tmp(74987) := x"0800";
    tmp(74988) := x"0800";
    tmp(74989) := x"2020";
    tmp(74990) := x"2020";
    tmp(74991) := x"2840";
    tmp(74992) := x"2040";
    tmp(74993) := x"0820";
    tmp(74994) := x"0020";
    tmp(74995) := x"0020";
    tmp(74996) := x"0020";
    tmp(74997) := x"0000";
    tmp(74998) := x"0000";
    tmp(74999) := x"0000";
    tmp(75000) := x"0000";
    tmp(75001) := x"0000";
    tmp(75002) := x"0000";
    tmp(75003) := x"0000";
    tmp(75004) := x"0000";
    tmp(75005) := x"0000";
    tmp(75006) := x"0000";
    tmp(75007) := x"0000";
    tmp(75008) := x"0000";
    tmp(75009) := x"0000";
    tmp(75010) := x"0000";
    tmp(75011) := x"0000";
    tmp(75012) := x"0020";
    tmp(75013) := x"0020";
    tmp(75014) := x"0020";
    tmp(75015) := x"0020";
    tmp(75016) := x"0020";
    tmp(75017) := x"0020";
    tmp(75018) := x"0020";
    tmp(75019) := x"0020";
    tmp(75020) := x"0020";
    tmp(75021) := x"0020";
    tmp(75022) := x"0020";
    tmp(75023) := x"0020";
    tmp(75024) := x"0020";
    tmp(75025) := x"0020";
    tmp(75026) := x"0020";
    tmp(75027) := x"0020";
    tmp(75028) := x"0020";
    tmp(75029) := x"0020";
    tmp(75030) := x"0020";
    tmp(75031) := x"0020";
    tmp(75032) := x"0020";
    tmp(75033) := x"0020";
    tmp(75034) := x"0020";
    tmp(75035) := x"0020";
    tmp(75036) := x"0020";
    tmp(75037) := x"0020";
    tmp(75038) := x"0020";
    tmp(75039) := x"0020";
    tmp(75040) := x"0020";
    tmp(75041) := x"0020";
    tmp(75042) := x"0020";
    tmp(75043) := x"0020";
    tmp(75044) := x"0000";
    tmp(75045) := x"0000";
    tmp(75046) := x"0000";
    tmp(75047) := x"0000";
    tmp(75048) := x"0000";
    tmp(75049) := x"0000";
    tmp(75050) := x"0000";
    tmp(75051) := x"0000";
    tmp(75052) := x"0000";
    tmp(75053) := x"0000";
    tmp(75054) := x"0000";
    tmp(75055) := x"0000";
    tmp(75056) := x"0000";
    tmp(75057) := x"0000";
    tmp(75058) := x"0000";
    tmp(75059) := x"0000";
    tmp(75060) := x"0000";
    tmp(75061) := x"0000";
    tmp(75062) := x"0000";
    tmp(75063) := x"0000";
    tmp(75064) := x"0000";
    tmp(75065) := x"0000";
    tmp(75066) := x"0000";
    tmp(75067) := x"0000";
    tmp(75068) := x"0000";
    tmp(75069) := x"0000";
    tmp(75070) := x"0000";
    tmp(75071) := x"0000";
    tmp(75072) := x"0000";
    tmp(75073) := x"0000";
    tmp(75074) := x"0000";
    tmp(75075) := x"0000";
    tmp(75076) := x"0000";
    tmp(75077) := x"0000";
    tmp(75078) := x"0000";
    tmp(75079) := x"0000";
    tmp(75080) := x"0000";
    tmp(75081) := x"0000";
    tmp(75082) := x"0000";
    tmp(75083) := x"0000";
    tmp(75084) := x"0000";
    tmp(75085) := x"0000";
    tmp(75086) := x"0000";
    tmp(75087) := x"0000";
    tmp(75088) := x"0000";
    tmp(75089) := x"0000";
    tmp(75090) := x"0000";
    tmp(75091) := x"0000";
    tmp(75092) := x"0000";
    tmp(75093) := x"0000";
    tmp(75094) := x"0000";
    tmp(75095) := x"0000";
    tmp(75096) := x"0000";
    tmp(75097) := x"0000";
    tmp(75098) := x"0000";
    tmp(75099) := x"0000";
    tmp(75100) := x"0000";
    tmp(75101) := x"0000";
    tmp(75102) := x"0000";
    tmp(75103) := x"0000";
    tmp(75104) := x"0000";
    tmp(75105) := x"0000";
    tmp(75106) := x"0000";
    tmp(75107) := x"0000";
    tmp(75108) := x"0000";
    tmp(75109) := x"0000";
    tmp(75110) := x"0000";
    tmp(75111) := x"0000";
    tmp(75112) := x"0000";
    tmp(75113) := x"0000";
    tmp(75114) := x"0000";
    tmp(75115) := x"0000";
    tmp(75116) := x"0000";
    tmp(75117) := x"0000";
    tmp(75118) := x"0000";
    tmp(75119) := x"0020";
    tmp(75120) := x"0000";
    tmp(75121) := x"0000";
    tmp(75122) := x"0000";
    tmp(75123) := x"0000";
    tmp(75124) := x"0000";
    tmp(75125) := x"0000";
    tmp(75126) := x"0000";
    tmp(75127) := x"0000";
    tmp(75128) := x"0000";
    tmp(75129) := x"0000";
    tmp(75130) := x"0000";
    tmp(75131) := x"0020";
    tmp(75132) := x"0020";
    tmp(75133) := x"0041";
    tmp(75134) := x"0041";
    tmp(75135) := x"0041";
    tmp(75136) := x"0040";
    tmp(75137) := x"0040";
    tmp(75138) := x"0020";
    tmp(75139) := x"0020";
    tmp(75140) := x"0020";
    tmp(75141) := x"0020";
    tmp(75142) := x"0020";
    tmp(75143) := x"0020";
    tmp(75144) := x"0020";
    tmp(75145) := x"0020";
    tmp(75146) := x"0020";
    tmp(75147) := x"0020";
    tmp(75148) := x"0020";
    tmp(75149) := x"0020";
    tmp(75150) := x"0020";
    tmp(75151) := x"0020";
    tmp(75152) := x"0040";
    tmp(75153) := x"0040";
    tmp(75154) := x"0040";
    tmp(75155) := x"0040";
    tmp(75156) := x"0040";
    tmp(75157) := x"0060";
    tmp(75158) := x"0060";
    tmp(75159) := x"0040";
    tmp(75160) := x"0040";
    tmp(75161) := x"0040";
    tmp(75162) := x"0040";
    tmp(75163) := x"0040";
    tmp(75164) := x"0060";
    tmp(75165) := x"0040";
    tmp(75166) := x"0040";
    tmp(75167) := x"0060";
    tmp(75168) := x"0060";
    tmp(75169) := x"0060";
    tmp(75170) := x"0060";
    tmp(75171) := x"0040";
    tmp(75172) := x"0040";
    tmp(75173) := x"0020";
    tmp(75174) := x"0020";
    tmp(75175) := x"0020";
    tmp(75176) := x"0020";
    tmp(75177) := x"0020";
    tmp(75178) := x"0020";
    tmp(75179) := x"0020";
    tmp(75180) := x"0020";
    tmp(75181) := x"0020";
    tmp(75182) := x"0020";
    tmp(75183) := x"0020";
    tmp(75184) := x"0020";
    tmp(75185) := x"0000";
    tmp(75186) := x"0000";
    tmp(75187) := x"0000";
    tmp(75188) := x"0000";
    tmp(75189) := x"0020";
    tmp(75190) := x"0820";
    tmp(75191) := x"0820";
    tmp(75192) := x"0820";
    tmp(75193) := x"0820";
    tmp(75194) := x"1000";
    tmp(75195) := x"1000";
    tmp(75196) := x"1000";
    tmp(75197) := x"1800";
    tmp(75198) := x"1800";
    tmp(75199) := x"1800";
    tmp(75200) := x"1800";
    tmp(75201) := x"1000";
    tmp(75202) := x"1800";
    tmp(75203) := x"1800";
    tmp(75204) := x"2000";
    tmp(75205) := x"2800";
    tmp(75206) := x"2800";
    tmp(75207) := x"2800";
    tmp(75208) := x"2800";
    tmp(75209) := x"2800";
    tmp(75210) := x"2800";
    tmp(75211) := x"2800";
    tmp(75212) := x"2800";
    tmp(75213) := x"2000";
    tmp(75214) := x"2000";
    tmp(75215) := x"2800";
    tmp(75216) := x"2800";
    tmp(75217) := x"2820";
    tmp(75218) := x"2820";
    tmp(75219) := x"2820";
    tmp(75220) := x"2020";
    tmp(75221) := x"1800";
    tmp(75222) := x"1000";
    tmp(75223) := x"0800";
    tmp(75224) := x"0800";
    tmp(75225) := x"1000";
    tmp(75226) := x"1800";
    tmp(75227) := x"2020";
    tmp(75228) := x"2820";
    tmp(75229) := x"3040";
    tmp(75230) := x"3040";
    tmp(75231) := x"1820";
    tmp(75232) := x"0820";
    tmp(75233) := x"0020";
    tmp(75234) := x"0020";
    tmp(75235) := x"0020";
    tmp(75236) := x"0000";
    tmp(75237) := x"0000";
    tmp(75238) := x"0000";
    tmp(75239) := x"0000";
    tmp(75240) := x"0000";
    tmp(75241) := x"0000";
    tmp(75242) := x"0000";
    tmp(75243) := x"0000";
    tmp(75244) := x"0000";
    tmp(75245) := x"0000";
    tmp(75246) := x"0000";
    tmp(75247) := x"0000";
    tmp(75248) := x"0000";
    tmp(75249) := x"0000";
    tmp(75250) := x"0000";
    tmp(75251) := x"0000";
    tmp(75252) := x"0000";
    tmp(75253) := x"0000";
    tmp(75254) := x"0000";
    tmp(75255) := x"0000";
    tmp(75256) := x"0000";
    tmp(75257) := x"0000";
    tmp(75258) := x"0020";
    tmp(75259) := x"0020";
    tmp(75260) := x"0020";
    tmp(75261) := x"0020";
    tmp(75262) := x"0020";
    tmp(75263) := x"0020";
    tmp(75264) := x"0020";
    tmp(75265) := x"0020";
    tmp(75266) := x"0020";
    tmp(75267) := x"0020";
    tmp(75268) := x"0020";
    tmp(75269) := x"0020";
    tmp(75270) := x"0020";
    tmp(75271) := x"0020";
    tmp(75272) := x"0020";
    tmp(75273) := x"0020";
    tmp(75274) := x"0020";
    tmp(75275) := x"0020";
    tmp(75276) := x"0020";
    tmp(75277) := x"0020";
    tmp(75278) := x"0020";
    tmp(75279) := x"0020";
    tmp(75280) := x"0000";
    tmp(75281) := x"0020";
    tmp(75282) := x"0000";
    tmp(75283) := x"0000";
    tmp(75284) := x"0000";
    tmp(75285) := x"0000";
    tmp(75286) := x"0000";
    tmp(75287) := x"0000";
    tmp(75288) := x"0000";
    tmp(75289) := x"0000";
    tmp(75290) := x"0000";
    tmp(75291) := x"0000";
    tmp(75292) := x"0000";
    tmp(75293) := x"0000";
    tmp(75294) := x"0000";
    tmp(75295) := x"0000";
    tmp(75296) := x"0000";
    tmp(75297) := x"0000";
    tmp(75298) := x"0000";
    tmp(75299) := x"0000";
    tmp(75300) := x"0000";
    tmp(75301) := x"0000";
    tmp(75302) := x"0000";
    tmp(75303) := x"0000";
    tmp(75304) := x"0000";
    tmp(75305) := x"0000";
    tmp(75306) := x"0000";
    tmp(75307) := x"0000";
    tmp(75308) := x"0000";
    tmp(75309) := x"0000";
    tmp(75310) := x"0000";
    tmp(75311) := x"0000";
    tmp(75312) := x"0000";
    tmp(75313) := x"0000";
    tmp(75314) := x"0000";
    tmp(75315) := x"0000";
    tmp(75316) := x"0000";
    tmp(75317) := x"0000";
    tmp(75318) := x"0000";
    tmp(75319) := x"0000";
    tmp(75320) := x"0000";
    tmp(75321) := x"0000";
    tmp(75322) := x"0000";
    tmp(75323) := x"0000";
    tmp(75324) := x"0000";
    tmp(75325) := x"0000";
    tmp(75326) := x"0000";
    tmp(75327) := x"0000";
    tmp(75328) := x"0000";
    tmp(75329) := x"0000";
    tmp(75330) := x"0000";
    tmp(75331) := x"0000";
    tmp(75332) := x"0000";
    tmp(75333) := x"0000";
    tmp(75334) := x"0000";
    tmp(75335) := x"0000";
    tmp(75336) := x"0000";
    tmp(75337) := x"0000";
    tmp(75338) := x"0000";
    tmp(75339) := x"0000";
    tmp(75340) := x"0000";
    tmp(75341) := x"0000";
    tmp(75342) := x"0000";
    tmp(75343) := x"0000";
    tmp(75344) := x"0000";
    tmp(75345) := x"0000";
    tmp(75346) := x"0000";
    tmp(75347) := x"0000";
    tmp(75348) := x"0000";
    tmp(75349) := x"0000";
    tmp(75350) := x"0000";
    tmp(75351) := x"0000";
    tmp(75352) := x"0000";
    tmp(75353) := x"0000";
    tmp(75354) := x"0000";
    tmp(75355) := x"0000";
    tmp(75356) := x"0000";
    tmp(75357) := x"0000";
    tmp(75358) := x"0000";
    tmp(75359) := x"0000";
    tmp(75360) := x"0000";
    tmp(75361) := x"0000";
    tmp(75362) := x"0000";
    tmp(75363) := x"0000";
    tmp(75364) := x"0000";
    tmp(75365) := x"0000";
    tmp(75366) := x"0000";
    tmp(75367) := x"0000";
    tmp(75368) := x"0000";
    tmp(75369) := x"0000";
    tmp(75370) := x"0000";
    tmp(75371) := x"0000";
    tmp(75372) := x"0000";
    tmp(75373) := x"0020";
    tmp(75374) := x"0020";
    tmp(75375) := x"0041";
    tmp(75376) := x"0041";
    tmp(75377) := x"0041";
    tmp(75378) := x"0040";
    tmp(75379) := x"0020";
    tmp(75380) := x"0020";
    tmp(75381) := x"0020";
    tmp(75382) := x"0020";
    tmp(75383) := x"0020";
    tmp(75384) := x"0020";
    tmp(75385) := x"0020";
    tmp(75386) := x"0020";
    tmp(75387) := x"0020";
    tmp(75388) := x"0020";
    tmp(75389) := x"0020";
    tmp(75390) := x"0020";
    tmp(75391) := x"0040";
    tmp(75392) := x"0040";
    tmp(75393) := x"0040";
    tmp(75394) := x"0040";
    tmp(75395) := x"0040";
    tmp(75396) := x"0040";
    tmp(75397) := x"0040";
    tmp(75398) := x"0040";
    tmp(75399) := x"0040";
    tmp(75400) := x"0040";
    tmp(75401) := x"0040";
    tmp(75402) := x"0020";
    tmp(75403) := x"0040";
    tmp(75404) := x"0040";
    tmp(75405) := x"0060";
    tmp(75406) := x"0860";
    tmp(75407) := x"0040";
    tmp(75408) := x"0060";
    tmp(75409) := x"0060";
    tmp(75410) := x"0040";
    tmp(75411) := x"0040";
    tmp(75412) := x"0020";
    tmp(75413) := x"0020";
    tmp(75414) := x"0020";
    tmp(75415) := x"0020";
    tmp(75416) := x"0020";
    tmp(75417) := x"0020";
    tmp(75418) := x"0020";
    tmp(75419) := x"0020";
    tmp(75420) := x"0020";
    tmp(75421) := x"0020";
    tmp(75422) := x"0820";
    tmp(75423) := x"0820";
    tmp(75424) := x"0820";
    tmp(75425) := x"0800";
    tmp(75426) := x"0800";
    tmp(75427) := x"0000";
    tmp(75428) := x"0000";
    tmp(75429) := x"0820";
    tmp(75430) := x"0800";
    tmp(75431) := x"0800";
    tmp(75432) := x"0800";
    tmp(75433) := x"1000";
    tmp(75434) := x"1000";
    tmp(75435) := x"1000";
    tmp(75436) := x"1000";
    tmp(75437) := x"1000";
    tmp(75438) := x"1000";
    tmp(75439) := x"1000";
    tmp(75440) := x"1000";
    tmp(75441) := x"1000";
    tmp(75442) := x"1000";
    tmp(75443) := x"1800";
    tmp(75444) := x"2000";
    tmp(75445) := x"2000";
    tmp(75446) := x"2800";
    tmp(75447) := x"2800";
    tmp(75448) := x"2800";
    tmp(75449) := x"2800";
    tmp(75450) := x"2800";
    tmp(75451) := x"2000";
    tmp(75452) := x"2000";
    tmp(75453) := x"1800";
    tmp(75454) := x"1800";
    tmp(75455) := x"2000";
    tmp(75456) := x"2000";
    tmp(75457) := x"2000";
    tmp(75458) := x"1800";
    tmp(75459) := x"1800";
    tmp(75460) := x"1800";
    tmp(75461) := x"1000";
    tmp(75462) := x"1000";
    tmp(75463) := x"1800";
    tmp(75464) := x"2020";
    tmp(75465) := x"2000";
    tmp(75466) := x"2000";
    tmp(75467) := x"3020";
    tmp(75468) := x"4040";
    tmp(75469) := x"2820";
    tmp(75470) := x"1020";
    tmp(75471) := x"0820";
    tmp(75472) := x"0020";
    tmp(75473) := x"0020";
    tmp(75474) := x"0020";
    tmp(75475) := x"0020";
    tmp(75476) := x"0020";
    tmp(75477) := x"0000";
    tmp(75478) := x"0000";
    tmp(75479) := x"0000";
    tmp(75480) := x"0000";
    tmp(75481) := x"0000";
    tmp(75482) := x"0000";
    tmp(75483) := x"0000";
    tmp(75484) := x"0000";
    tmp(75485) := x"0000";
    tmp(75486) := x"0000";
    tmp(75487) := x"0000";
    tmp(75488) := x"0000";
    tmp(75489) := x"0000";
    tmp(75490) := x"0000";
    tmp(75491) := x"0000";
    tmp(75492) := x"0000";
    tmp(75493) := x"0000";
    tmp(75494) := x"0000";
    tmp(75495) := x"0000";
    tmp(75496) := x"0000";
    tmp(75497) := x"0000";
    tmp(75498) := x"0000";
    tmp(75499) := x"0000";
    tmp(75500) := x"0000";
    tmp(75501) := x"0000";
    tmp(75502) := x"0000";
    tmp(75503) := x"0000";
    tmp(75504) := x"0000";
    tmp(75505) := x"0000";
    tmp(75506) := x"0000";
    tmp(75507) := x"0020";
    tmp(75508) := x"0000";
    tmp(75509) := x"0000";
    tmp(75510) := x"0020";
    tmp(75511) := x"0000";
    tmp(75512) := x"0000";
    tmp(75513) := x"0000";
    tmp(75514) := x"0000";
    tmp(75515) := x"0000";
    tmp(75516) := x"0000";
    tmp(75517) := x"0000";
    tmp(75518) := x"0000";
    tmp(75519) := x"0020";
    tmp(75520) := x"0000";
    tmp(75521) := x"0000";
    tmp(75522) := x"0000";
    tmp(75523) := x"0000";
    tmp(75524) := x"0000";
    tmp(75525) := x"0000";
    tmp(75526) := x"0000";
    tmp(75527) := x"0000";
    tmp(75528) := x"0000";
    tmp(75529) := x"0000";
    tmp(75530) := x"0000";
    tmp(75531) := x"0000";
    tmp(75532) := x"0000";
    tmp(75533) := x"0000";
    tmp(75534) := x"0000";
    tmp(75535) := x"0000";
    tmp(75536) := x"0000";
    tmp(75537) := x"0000";
    tmp(75538) := x"0000";
    tmp(75539) := x"0000";
    tmp(75540) := x"0000";
    tmp(75541) := x"0000";
    tmp(75542) := x"0000";
    tmp(75543) := x"0000";
    tmp(75544) := x"0000";
    tmp(75545) := x"0000";
    tmp(75546) := x"0000";
    tmp(75547) := x"0000";
    tmp(75548) := x"0000";
    tmp(75549) := x"0000";
    tmp(75550) := x"0000";
    tmp(75551) := x"0000";
    tmp(75552) := x"0000";
    tmp(75553) := x"0000";
    tmp(75554) := x"0000";
    tmp(75555) := x"0000";
    tmp(75556) := x"0000";
    tmp(75557) := x"0000";
    tmp(75558) := x"0000";
    tmp(75559) := x"0000";
    tmp(75560) := x"0000";
    tmp(75561) := x"0000";
    tmp(75562) := x"0000";
    tmp(75563) := x"0000";
    tmp(75564) := x"0000";
    tmp(75565) := x"0000";
    tmp(75566) := x"0000";
    tmp(75567) := x"0000";
    tmp(75568) := x"0000";
    tmp(75569) := x"0000";
    tmp(75570) := x"0000";
    tmp(75571) := x"0000";
    tmp(75572) := x"0000";
    tmp(75573) := x"0000";
    tmp(75574) := x"0000";
    tmp(75575) := x"0000";
    tmp(75576) := x"0000";
    tmp(75577) := x"0000";
    tmp(75578) := x"0000";
    tmp(75579) := x"0000";
    tmp(75580) := x"0000";
    tmp(75581) := x"0000";
    tmp(75582) := x"0000";
    tmp(75583) := x"0000";
    tmp(75584) := x"0000";
    tmp(75585) := x"0000";
    tmp(75586) := x"0000";
    tmp(75587) := x"0000";
    tmp(75588) := x"0000";
    tmp(75589) := x"0000";
    tmp(75590) := x"0000";
    tmp(75591) := x"0000";
    tmp(75592) := x"0000";
    tmp(75593) := x"0000";
    tmp(75594) := x"0000";
    tmp(75595) := x"0000";
    tmp(75596) := x"0000";
    tmp(75597) := x"0000";
    tmp(75598) := x"0000";
    tmp(75599) := x"0000";
    tmp(75600) := x"0000";
    tmp(75601) := x"0000";
    tmp(75602) := x"0000";
    tmp(75603) := x"0000";
    tmp(75604) := x"0000";
    tmp(75605) := x"0000";
    tmp(75606) := x"0000";
    tmp(75607) := x"0000";
    tmp(75608) := x"0000";
    tmp(75609) := x"0000";
    tmp(75610) := x"0000";
    tmp(75611) := x"0000";
    tmp(75612) := x"0000";
    tmp(75613) := x"0000";
    tmp(75614) := x"0000";
    tmp(75615) := x"0020";
    tmp(75616) := x"0020";
    tmp(75617) := x"0040";
    tmp(75618) := x"0040";
    tmp(75619) := x"0040";
    tmp(75620) := x"0020";
    tmp(75621) := x"0020";
    tmp(75622) := x"0020";
    tmp(75623) := x"0020";
    tmp(75624) := x"0020";
    tmp(75625) := x"0020";
    tmp(75626) := x"0020";
    tmp(75627) := x"0020";
    tmp(75628) := x"0020";
    tmp(75629) := x"0020";
    tmp(75630) := x"0040";
    tmp(75631) := x"0040";
    tmp(75632) := x"0040";
    tmp(75633) := x"0040";
    tmp(75634) := x"0040";
    tmp(75635) := x"0040";
    tmp(75636) := x"0040";
    tmp(75637) := x"0040";
    tmp(75638) := x"0040";
    tmp(75639) := x"0040";
    tmp(75640) := x"0040";
    tmp(75641) := x"0020";
    tmp(75642) := x"0020";
    tmp(75643) := x"0040";
    tmp(75644) := x"0020";
    tmp(75645) := x"0020";
    tmp(75646) := x"0040";
    tmp(75647) := x"0040";
    tmp(75648) := x"0040";
    tmp(75649) := x"0040";
    tmp(75650) := x"0040";
    tmp(75651) := x"0040";
    tmp(75652) := x"0040";
    tmp(75653) := x"0040";
    tmp(75654) := x"0820";
    tmp(75655) := x"0820";
    tmp(75656) := x"0800";
    tmp(75657) := x"0800";
    tmp(75658) := x"0800";
    tmp(75659) := x"0800";
    tmp(75660) := x"0000";
    tmp(75661) := x"0000";
    tmp(75662) := x"0820";
    tmp(75663) := x"0820";
    tmp(75664) := x"0820";
    tmp(75665) := x"0800";
    tmp(75666) := x"0800";
    tmp(75667) := x"0800";
    tmp(75668) := x"0800";
    tmp(75669) := x"0800";
    tmp(75670) := x"0800";
    tmp(75671) := x"0800";
    tmp(75672) := x"0800";
    tmp(75673) := x"1000";
    tmp(75674) := x"1000";
    tmp(75675) := x"1000";
    tmp(75676) := x"0800";
    tmp(75677) := x"1000";
    tmp(75678) := x"1000";
    tmp(75679) := x"1000";
    tmp(75680) := x"1000";
    tmp(75681) := x"1000";
    tmp(75682) := x"1000";
    tmp(75683) := x"1800";
    tmp(75684) := x"1800";
    tmp(75685) := x"2000";
    tmp(75686) := x"2800";
    tmp(75687) := x"2000";
    tmp(75688) := x"2000";
    tmp(75689) := x"2000";
    tmp(75690) := x"2000";
    tmp(75691) := x"2000";
    tmp(75692) := x"1800";
    tmp(75693) := x"1800";
    tmp(75694) := x"1800";
    tmp(75695) := x"2000";
    tmp(75696) := x"2000";
    tmp(75697) := x"2000";
    tmp(75698) := x"2000";
    tmp(75699) := x"2800";
    tmp(75700) := x"2000";
    tmp(75701) := x"2000";
    tmp(75702) := x"2000";
    tmp(75703) := x"2820";
    tmp(75704) := x"2000";
    tmp(75705) := x"1800";
    tmp(75706) := x"2820";
    tmp(75707) := x"3840";
    tmp(75708) := x"3020";
    tmp(75709) := x"1020";
    tmp(75710) := x"0820";
    tmp(75711) := x"0020";
    tmp(75712) := x"0020";
    tmp(75713) := x"0020";
    tmp(75714) := x"0020";
    tmp(75715) := x"0020";
    tmp(75716) := x"0000";
    tmp(75717) := x"0000";
    tmp(75718) := x"0000";
    tmp(75719) := x"0000";
    tmp(75720) := x"0000";
    tmp(75721) := x"0000";
    tmp(75722) := x"0000";
    tmp(75723) := x"0000";
    tmp(75724) := x"0000";
    tmp(75725) := x"0000";
    tmp(75726) := x"0000";
    tmp(75727) := x"0000";
    tmp(75728) := x"0000";
    tmp(75729) := x"0000";
    tmp(75730) := x"0000";
    tmp(75731) := x"0000";
    tmp(75732) := x"0000";
    tmp(75733) := x"0000";
    tmp(75734) := x"0000";
    tmp(75735) := x"0000";
    tmp(75736) := x"0000";
    tmp(75737) := x"0000";
    tmp(75738) := x"0000";
    tmp(75739) := x"0000";
    tmp(75740) := x"0000";
    tmp(75741) := x"0000";
    tmp(75742) := x"0000";
    tmp(75743) := x"0000";
    tmp(75744) := x"0000";
    tmp(75745) := x"0000";
    tmp(75746) := x"0000";
    tmp(75747) := x"0000";
    tmp(75748) := x"0000";
    tmp(75749) := x"0000";
    tmp(75750) := x"0000";
    tmp(75751) := x"0000";
    tmp(75752) := x"0000";
    tmp(75753) := x"0000";
    tmp(75754) := x"0000";
    tmp(75755) := x"0000";
    tmp(75756) := x"0000";
    tmp(75757) := x"0000";
    tmp(75758) := x"0000";
    tmp(75759) := x"0000";
    tmp(75760) := x"0000";
    tmp(75761) := x"0000";
    tmp(75762) := x"0000";
    tmp(75763) := x"0000";
    tmp(75764) := x"0000";
    tmp(75765) := x"0000";
    tmp(75766) := x"0000";
    tmp(75767) := x"0000";
    tmp(75768) := x"0000";
    tmp(75769) := x"0000";
    tmp(75770) := x"0000";
    tmp(75771) := x"0000";
    tmp(75772) := x"0000";
    tmp(75773) := x"0000";
    tmp(75774) := x"0000";
    tmp(75775) := x"0000";
    tmp(75776) := x"0000";
    tmp(75777) := x"0000";
    tmp(75778) := x"0000";
    tmp(75779) := x"0000";
    tmp(75780) := x"0000";
    tmp(75781) := x"0000";
    tmp(75782) := x"0000";
    tmp(75783) := x"0000";
    tmp(75784) := x"0000";
    tmp(75785) := x"0000";
    tmp(75786) := x"0000";
    tmp(75787) := x"0000";
    tmp(75788) := x"0000";
    tmp(75789) := x"0000";
    tmp(75790) := x"0000";
    tmp(75791) := x"0000";
    tmp(75792) := x"0000";
    tmp(75793) := x"0000";
    tmp(75794) := x"0000";
    tmp(75795) := x"0000";
    tmp(75796) := x"0000";
    tmp(75797) := x"0000";
    tmp(75798) := x"0000";
    tmp(75799) := x"0000";
    tmp(75800) := x"0000";
    tmp(75801) := x"0000";
    tmp(75802) := x"0000";
    tmp(75803) := x"0000";
    tmp(75804) := x"0000";
    tmp(75805) := x"0000";
    tmp(75806) := x"0000";
    tmp(75807) := x"0000";
    tmp(75808) := x"0000";
    tmp(75809) := x"0000";
    tmp(75810) := x"0000";
    tmp(75811) := x"0000";
    tmp(75812) := x"0000";
    tmp(75813) := x"0000";
    tmp(75814) := x"0000";
    tmp(75815) := x"0000";
    tmp(75816) := x"0000";
    tmp(75817) := x"0000";
    tmp(75818) := x"0000";
    tmp(75819) := x"0000";
    tmp(75820) := x"0000";
    tmp(75821) := x"0000";
    tmp(75822) := x"0000";
    tmp(75823) := x"0000";
    tmp(75824) := x"0000";
    tmp(75825) := x"0000";
    tmp(75826) := x"0000";
    tmp(75827) := x"0000";
    tmp(75828) := x"0000";
    tmp(75829) := x"0000";
    tmp(75830) := x"0000";
    tmp(75831) := x"0000";
    tmp(75832) := x"0000";
    tmp(75833) := x"0000";
    tmp(75834) := x"0000";
    tmp(75835) := x"0000";
    tmp(75836) := x"0000";
    tmp(75837) := x"0000";
    tmp(75838) := x"0000";
    tmp(75839) := x"0000";
    tmp(75840) := x"0000";
    tmp(75841) := x"0000";
    tmp(75842) := x"0000";
    tmp(75843) := x"0000";
    tmp(75844) := x"0000";
    tmp(75845) := x"0020";
    tmp(75846) := x"0020";
    tmp(75847) := x"0020";
    tmp(75848) := x"0020";
    tmp(75849) := x"0020";
    tmp(75850) := x"0020";
    tmp(75851) := x"0020";
    tmp(75852) := x"0000";
    tmp(75853) := x"0000";
    tmp(75854) := x"0000";
    tmp(75855) := x"0000";
    tmp(75856) := x"0000";
    tmp(75857) := x"0020";
    tmp(75858) := x"0020";
    tmp(75859) := x"0020";
    tmp(75860) := x"0020";
    tmp(75861) := x"0040";
    tmp(75862) := x"0020";
    tmp(75863) := x"0020";
    tmp(75864) := x"0020";
    tmp(75865) := x"0020";
    tmp(75866) := x"0020";
    tmp(75867) := x"0020";
    tmp(75868) := x"0020";
    tmp(75869) := x"0020";
    tmp(75870) := x"0020";
    tmp(75871) := x"0020";
    tmp(75872) := x"0040";
    tmp(75873) := x"0040";
    tmp(75874) := x"0040";
    tmp(75875) := x"0040";
    tmp(75876) := x"0040";
    tmp(75877) := x"0040";
    tmp(75878) := x"0040";
    tmp(75879) := x"0040";
    tmp(75880) := x"0040";
    tmp(75881) := x"0020";
    tmp(75882) := x"0040";
    tmp(75883) := x"0040";
    tmp(75884) := x"0020";
    tmp(75885) := x"0020";
    tmp(75886) := x"0020";
    tmp(75887) := x"0020";
    tmp(75888) := x"0040";
    tmp(75889) := x"0040";
    tmp(75890) := x"0040";
    tmp(75891) := x"0840";
    tmp(75892) := x"0840";
    tmp(75893) := x"0840";
    tmp(75894) := x"0840";
    tmp(75895) := x"0820";
    tmp(75896) := x"0800";
    tmp(75897) := x"0800";
    tmp(75898) := x"0800";
    tmp(75899) := x"0800";
    tmp(75900) := x"0800";
    tmp(75901) := x"0820";
    tmp(75902) := x"0820";
    tmp(75903) := x"0820";
    tmp(75904) := x"0820";
    tmp(75905) := x"0820";
    tmp(75906) := x"0820";
    tmp(75907) := x"0820";
    tmp(75908) := x"0800";
    tmp(75909) := x"0800";
    tmp(75910) := x"0800";
    tmp(75911) := x"0800";
    tmp(75912) := x"1000";
    tmp(75913) := x"1000";
    tmp(75914) := x"1000";
    tmp(75915) := x"0800";
    tmp(75916) := x"0800";
    tmp(75917) := x"1000";
    tmp(75918) := x"1000";
    tmp(75919) := x"1000";
    tmp(75920) := x"1800";
    tmp(75921) := x"1800";
    tmp(75922) := x"1000";
    tmp(75923) := x"1000";
    tmp(75924) := x"1000";
    tmp(75925) := x"1800";
    tmp(75926) := x"2000";
    tmp(75927) := x"2000";
    tmp(75928) := x"2800";
    tmp(75929) := x"2800";
    tmp(75930) := x"2820";
    tmp(75931) := x"2820";
    tmp(75932) := x"2820";
    tmp(75933) := x"2820";
    tmp(75934) := x"3020";
    tmp(75935) := x"3020";
    tmp(75936) := x"3820";
    tmp(75937) := x"3820";
    tmp(75938) := x"3020";
    tmp(75939) := x"2000";
    tmp(75940) := x"1800";
    tmp(75941) := x"2000";
    tmp(75942) := x"2820";
    tmp(75943) := x"2800";
    tmp(75944) := x"1000";
    tmp(75945) := x"2000";
    tmp(75946) := x"3020";
    tmp(75947) := x"2020";
    tmp(75948) := x"1000";
    tmp(75949) := x"0820";
    tmp(75950) := x"0020";
    tmp(75951) := x"0020";
    tmp(75952) := x"0020";
    tmp(75953) := x"0020";
    tmp(75954) := x"0020";
    tmp(75955) := x"0020";
    tmp(75956) := x"0000";
    tmp(75957) := x"0000";
    tmp(75958) := x"0000";
    tmp(75959) := x"0000";
    tmp(75960) := x"0000";
    tmp(75961) := x"0000";
    tmp(75962) := x"0000";
    tmp(75963) := x"0000";
    tmp(75964) := x"0000";
    tmp(75965) := x"0000";
    tmp(75966) := x"0000";
    tmp(75967) := x"0000";
    tmp(75968) := x"0000";
    tmp(75969) := x"0000";
    tmp(75970) := x"0000";
    tmp(75971) := x"0000";
    tmp(75972) := x"0000";
    tmp(75973) := x"0000";
    tmp(75974) := x"0000";
    tmp(75975) := x"0000";
    tmp(75976) := x"0000";
    tmp(75977) := x"0000";
    tmp(75978) := x"0000";
    tmp(75979) := x"0000";
    tmp(75980) := x"0000";
    tmp(75981) := x"0000";
    tmp(75982) := x"0000";
    tmp(75983) := x"0000";
    tmp(75984) := x"0000";
    tmp(75985) := x"0000";
    tmp(75986) := x"0000";
    tmp(75987) := x"0000";
    tmp(75988) := x"0000";
    tmp(75989) := x"0000";
    tmp(75990) := x"0000";
    tmp(75991) := x"0000";
    tmp(75992) := x"0000";
    tmp(75993) := x"0000";
    tmp(75994) := x"0000";
    tmp(75995) := x"0000";
    tmp(75996) := x"0000";
    tmp(75997) := x"0000";
    tmp(75998) := x"0000";
    tmp(75999) := x"0000";
    tmp(76000) := x"0000";
    tmp(76001) := x"0000";
    tmp(76002) := x"0000";
    tmp(76003) := x"0000";
    tmp(76004) := x"0000";
    tmp(76005) := x"0000";
    tmp(76006) := x"0000";
    tmp(76007) := x"0000";
    tmp(76008) := x"0000";
    tmp(76009) := x"0000";
    tmp(76010) := x"0000";
    tmp(76011) := x"0000";
    tmp(76012) := x"0000";
    tmp(76013) := x"0000";
    tmp(76014) := x"0000";
    tmp(76015) := x"0000";
    tmp(76016) := x"0000";
    tmp(76017) := x"0000";
    tmp(76018) := x"0000";
    tmp(76019) := x"0000";
    tmp(76020) := x"0000";
    tmp(76021) := x"0000";
    tmp(76022) := x"0000";
    tmp(76023) := x"0000";
    tmp(76024) := x"0000";
    tmp(76025) := x"0000";
    tmp(76026) := x"0000";
    tmp(76027) := x"0000";
    tmp(76028) := x"0000";
    tmp(76029) := x"0000";
    tmp(76030) := x"0000";
    tmp(76031) := x"0000";
    tmp(76032) := x"0000";
    tmp(76033) := x"0000";
    tmp(76034) := x"0000";
    tmp(76035) := x"0000";
    tmp(76036) := x"0000";
    tmp(76037) := x"0000";
    tmp(76038) := x"0000";
    tmp(76039) := x"0000";
    tmp(76040) := x"0000";
    tmp(76041) := x"0000";
    tmp(76042) := x"0000";
    tmp(76043) := x"0000";
    tmp(76044) := x"0000";
    tmp(76045) := x"0000";
    tmp(76046) := x"0000";
    tmp(76047) := x"0000";
    tmp(76048) := x"0000";
    tmp(76049) := x"0000";
    tmp(76050) := x"0000";
    tmp(76051) := x"0000";
    tmp(76052) := x"0000";
    tmp(76053) := x"0000";
    tmp(76054) := x"0000";
    tmp(76055) := x"0000";
    tmp(76056) := x"0000";
    tmp(76057) := x"0000";
    tmp(76058) := x"0000";
    tmp(76059) := x"0000";
    tmp(76060) := x"0000";
    tmp(76061) := x"0000";
    tmp(76062) := x"0000";
    tmp(76063) := x"0000";
    tmp(76064) := x"0000";
    tmp(76065) := x"0000";
    tmp(76066) := x"0000";
    tmp(76067) := x"0000";
    tmp(76068) := x"0000";
    tmp(76069) := x"0000";
    tmp(76070) := x"0000";
    tmp(76071) := x"0000";
    tmp(76072) := x"0000";
    tmp(76073) := x"0000";
    tmp(76074) := x"0000";
    tmp(76075) := x"0000";
    tmp(76076) := x"0000";
    tmp(76077) := x"0000";
    tmp(76078) := x"0000";
    tmp(76079) := x"0000";
    tmp(76080) := x"0000";
    tmp(76081) := x"0000";
    tmp(76082) := x"0000";
    tmp(76083) := x"0000";
    tmp(76084) := x"0020";
    tmp(76085) := x"0020";
    tmp(76086) := x"0021";
    tmp(76087) := x"0041";
    tmp(76088) := x"0041";
    tmp(76089) := x"0041";
    tmp(76090) := x"0041";
    tmp(76091) := x"0041";
    tmp(76092) := x"0040";
    tmp(76093) := x"0020";
    tmp(76094) := x"0020";
    tmp(76095) := x"0020";
    tmp(76096) := x"0020";
    tmp(76097) := x"0020";
    tmp(76098) := x"0020";
    tmp(76099) := x"0020";
    tmp(76100) := x"0020";
    tmp(76101) := x"0020";
    tmp(76102) := x"0040";
    tmp(76103) := x"0040";
    tmp(76104) := x"0020";
    tmp(76105) := x"0020";
    tmp(76106) := x"0020";
    tmp(76107) := x"0020";
    tmp(76108) := x"0020";
    tmp(76109) := x"0020";
    tmp(76110) := x"0020";
    tmp(76111) := x"0020";
    tmp(76112) := x"0020";
    tmp(76113) := x"0020";
    tmp(76114) := x"0020";
    tmp(76115) := x"0020";
    tmp(76116) := x"0040";
    tmp(76117) := x"0040";
    tmp(76118) := x"0040";
    tmp(76119) := x"0040";
    tmp(76120) := x"0040";
    tmp(76121) := x"0040";
    tmp(76122) := x"0040";
    tmp(76123) := x"0040";
    tmp(76124) := x"0840";
    tmp(76125) := x"0040";
    tmp(76126) := x"0040";
    tmp(76127) := x"0040";
    tmp(76128) := x"0040";
    tmp(76129) := x"0040";
    tmp(76130) := x"0040";
    tmp(76131) := x"0040";
    tmp(76132) := x"0840";
    tmp(76133) := x"0840";
    tmp(76134) := x"0840";
    tmp(76135) := x"0840";
    tmp(76136) := x"0820";
    tmp(76137) := x"0800";
    tmp(76138) := x"0800";
    tmp(76139) := x"0800";
    tmp(76140) := x"0820";
    tmp(76141) := x"0820";
    tmp(76142) := x"0820";
    tmp(76143) := x"0820";
    tmp(76144) := x"0820";
    tmp(76145) := x"0820";
    tmp(76146) := x"0820";
    tmp(76147) := x"1020";
    tmp(76148) := x"1020";
    tmp(76149) := x"0800";
    tmp(76150) := x"0800";
    tmp(76151) := x"1000";
    tmp(76152) := x"1000";
    tmp(76153) := x"1000";
    tmp(76154) := x"0800";
    tmp(76155) := x"1000";
    tmp(76156) := x"1000";
    tmp(76157) := x"1000";
    tmp(76158) := x"1000";
    tmp(76159) := x"1000";
    tmp(76160) := x"1800";
    tmp(76161) := x"1000";
    tmp(76162) := x"1000";
    tmp(76163) := x"1000";
    tmp(76164) := x"1000";
    tmp(76165) := x"1800";
    tmp(76166) := x"2020";
    tmp(76167) := x"2820";
    tmp(76168) := x"2820";
    tmp(76169) := x"2820";
    tmp(76170) := x"2820";
    tmp(76171) := x"2000";
    tmp(76172) := x"2000";
    tmp(76173) := x"2820";
    tmp(76174) := x"2820";
    tmp(76175) := x"2820";
    tmp(76176) := x"2820";
    tmp(76177) := x"2000";
    tmp(76178) := x"1000";
    tmp(76179) := x"1000";
    tmp(76180) := x"2000";
    tmp(76181) := x"3020";
    tmp(76182) := x"3020";
    tmp(76183) := x"1800";
    tmp(76184) := x"1000";
    tmp(76185) := x"2020";
    tmp(76186) := x"1800";
    tmp(76187) := x"1000";
    tmp(76188) := x"1000";
    tmp(76189) := x"0820";
    tmp(76190) := x"0020";
    tmp(76191) := x"0020";
    tmp(76192) := x"0020";
    tmp(76193) := x"0020";
    tmp(76194) := x"0020";
    tmp(76195) := x"0020";
    tmp(76196) := x"0020";
    tmp(76197) := x"0000";
    tmp(76198) := x"0000";
    tmp(76199) := x"0000";
    tmp(76200) := x"0000";
    tmp(76201) := x"0000";
    tmp(76202) := x"0000";
    tmp(76203) := x"0000";
    tmp(76204) := x"0000";
    tmp(76205) := x"0000";
    tmp(76206) := x"0000";
    tmp(76207) := x"0000";
    tmp(76208) := x"0000";
    tmp(76209) := x"0000";
    tmp(76210) := x"0000";
    tmp(76211) := x"0000";
    tmp(76212) := x"0000";
    tmp(76213) := x"0000";
    tmp(76214) := x"0000";
    tmp(76215) := x"0000";
    tmp(76216) := x"0000";
    tmp(76217) := x"0000";
    tmp(76218) := x"0000";
    tmp(76219) := x"0000";
    tmp(76220) := x"0000";
    tmp(76221) := x"0000";
    tmp(76222) := x"0000";
    tmp(76223) := x"0000";
    tmp(76224) := x"0000";
    tmp(76225) := x"0000";
    tmp(76226) := x"0000";
    tmp(76227) := x"0000";
    tmp(76228) := x"0000";
    tmp(76229) := x"0000";
    tmp(76230) := x"0000";
    tmp(76231) := x"0000";
    tmp(76232) := x"0000";
    tmp(76233) := x"0000";
    tmp(76234) := x"0000";
    tmp(76235) := x"0000";
    tmp(76236) := x"0000";
    tmp(76237) := x"0000";
    tmp(76238) := x"0000";
    tmp(76239) := x"0000";
    tmp(76240) := x"0000";
    tmp(76241) := x"0000";
    tmp(76242) := x"0000";
    tmp(76243) := x"0000";
    tmp(76244) := x"0000";
    tmp(76245) := x"0000";
    tmp(76246) := x"0000";
    tmp(76247) := x"0000";
    tmp(76248) := x"0000";
    tmp(76249) := x"0000";
    tmp(76250) := x"0000";
    tmp(76251) := x"0000";
    tmp(76252) := x"0000";
    tmp(76253) := x"0000";
    tmp(76254) := x"0000";
    tmp(76255) := x"0000";
    tmp(76256) := x"0000";
    tmp(76257) := x"0000";
    tmp(76258) := x"0000";
    tmp(76259) := x"0000";
    tmp(76260) := x"0000";
    tmp(76261) := x"0000";
    tmp(76262) := x"0000";
    tmp(76263) := x"0000";
    tmp(76264) := x"0000";
    tmp(76265) := x"0000";
    tmp(76266) := x"0000";
    tmp(76267) := x"0000";
    tmp(76268) := x"0000";
    tmp(76269) := x"0000";
    tmp(76270) := x"0000";
    tmp(76271) := x"0000";
    tmp(76272) := x"0000";
    tmp(76273) := x"0000";
    tmp(76274) := x"0000";
    tmp(76275) := x"0000";
    tmp(76276) := x"0000";
    tmp(76277) := x"0000";
    tmp(76278) := x"0000";
    tmp(76279) := x"0000";
    tmp(76280) := x"0000";
    tmp(76281) := x"0000";
    tmp(76282) := x"0000";
    tmp(76283) := x"0000";
    tmp(76284) := x"0000";
    tmp(76285) := x"0000";
    tmp(76286) := x"0000";
    tmp(76287) := x"0000";
    tmp(76288) := x"0000";
    tmp(76289) := x"0000";
    tmp(76290) := x"0000";
    tmp(76291) := x"0000";
    tmp(76292) := x"0000";
    tmp(76293) := x"0000";
    tmp(76294) := x"0000";
    tmp(76295) := x"0000";
    tmp(76296) := x"0000";
    tmp(76297) := x"0000";
    tmp(76298) := x"0000";
    tmp(76299) := x"0000";
    tmp(76300) := x"0000";
    tmp(76301) := x"0000";
    tmp(76302) := x"0000";
    tmp(76303) := x"0000";
    tmp(76304) := x"0000";
    tmp(76305) := x"0000";
    tmp(76306) := x"0000";
    tmp(76307) := x"0000";
    tmp(76308) := x"0000";
    tmp(76309) := x"0000";
    tmp(76310) := x"0000";
    tmp(76311) := x"0000";
    tmp(76312) := x"0000";
    tmp(76313) := x"0000";
    tmp(76314) := x"0000";
    tmp(76315) := x"0000";
    tmp(76316) := x"0000";
    tmp(76317) := x"0000";
    tmp(76318) := x"0000";
    tmp(76319) := x"0000";
    tmp(76320) := x"0000";
    tmp(76321) := x"0000";
    tmp(76322) := x"0000";
    tmp(76323) := x"0000";
    tmp(76324) := x"0020";
    tmp(76325) := x"0020";
    tmp(76326) := x"0020";
    tmp(76327) := x"0041";
    tmp(76328) := x"0041";
    tmp(76329) := x"0041";
    tmp(76330) := x"0041";
    tmp(76331) := x"0040";
    tmp(76332) := x"0040";
    tmp(76333) := x"0040";
    tmp(76334) := x"0040";
    tmp(76335) := x"0040";
    tmp(76336) := x"0040";
    tmp(76337) := x"0040";
    tmp(76338) := x"0040";
    tmp(76339) := x"0020";
    tmp(76340) := x"0020";
    tmp(76341) := x"0020";
    tmp(76342) := x"0040";
    tmp(76343) := x"0040";
    tmp(76344) := x"0040";
    tmp(76345) := x"0020";
    tmp(76346) := x"0020";
    tmp(76347) := x"0020";
    tmp(76348) := x"0020";
    tmp(76349) := x"0020";
    tmp(76350) := x"0020";
    tmp(76351) := x"0020";
    tmp(76352) := x"0020";
    tmp(76353) := x"0020";
    tmp(76354) := x"0020";
    tmp(76355) := x"0040";
    tmp(76356) := x"0020";
    tmp(76357) := x"0020";
    tmp(76358) := x"0020";
    tmp(76359) := x"0020";
    tmp(76360) := x"0020";
    tmp(76361) := x"0020";
    tmp(76362) := x"0020";
    tmp(76363) := x"0020";
    tmp(76364) := x"0040";
    tmp(76365) := x"0840";
    tmp(76366) := x"0840";
    tmp(76367) := x"0040";
    tmp(76368) := x"0040";
    tmp(76369) := x"0040";
    tmp(76370) := x"0040";
    tmp(76371) := x"0040";
    tmp(76372) := x"0040";
    tmp(76373) := x"0040";
    tmp(76374) := x"0040";
    tmp(76375) := x"0040";
    tmp(76376) := x"0840";
    tmp(76377) := x"0820";
    tmp(76378) := x"0820";
    tmp(76379) := x"0820";
    tmp(76380) := x"0820";
    tmp(76381) := x"0820";
    tmp(76382) := x"0820";
    tmp(76383) := x"0820";
    tmp(76384) := x"0820";
    tmp(76385) := x"1020";
    tmp(76386) := x"1020";
    tmp(76387) := x"1020";
    tmp(76388) := x"1020";
    tmp(76389) := x"1020";
    tmp(76390) := x"1000";
    tmp(76391) := x"1000";
    tmp(76392) := x"1000";
    tmp(76393) := x"1000";
    tmp(76394) := x"1000";
    tmp(76395) := x"1000";
    tmp(76396) := x"1000";
    tmp(76397) := x"1000";
    tmp(76398) := x"1000";
    tmp(76399) := x"1000";
    tmp(76400) := x"1000";
    tmp(76401) := x"1000";
    tmp(76402) := x"1000";
    tmp(76403) := x"1000";
    tmp(76404) := x"1800";
    tmp(76405) := x"2020";
    tmp(76406) := x"2820";
    tmp(76407) := x"2820";
    tmp(76408) := x"2820";
    tmp(76409) := x"2000";
    tmp(76410) := x"1800";
    tmp(76411) := x"1800";
    tmp(76412) := x"2000";
    tmp(76413) := x"2800";
    tmp(76414) := x"2000";
    tmp(76415) := x"2000";
    tmp(76416) := x"2000";
    tmp(76417) := x"1800";
    tmp(76418) := x"1000";
    tmp(76419) := x"1800";
    tmp(76420) := x"2820";
    tmp(76421) := x"2820";
    tmp(76422) := x"1000";
    tmp(76423) := x"0800";
    tmp(76424) := x"1000";
    tmp(76425) := x"1000";
    tmp(76426) := x"1000";
    tmp(76427) := x"1000";
    tmp(76428) := x"1020";
    tmp(76429) := x"0820";
    tmp(76430) := x"0020";
    tmp(76431) := x"0020";
    tmp(76432) := x"0020";
    tmp(76433) := x"0020";
    tmp(76434) := x"0020";
    tmp(76435) := x"0020";
    tmp(76436) := x"0000";
    tmp(76437) := x"0000";
    tmp(76438) := x"0000";
    tmp(76439) := x"0000";
    tmp(76440) := x"0000";
    tmp(76441) := x"0000";
    tmp(76442) := x"0000";
    tmp(76443) := x"0000";
    tmp(76444) := x"0000";
    tmp(76445) := x"0000";
    tmp(76446) := x"0000";
    tmp(76447) := x"0000";
    tmp(76448) := x"0000";
    tmp(76449) := x"0000";
    tmp(76450) := x"0000";
    tmp(76451) := x"0000";
    tmp(76452) := x"0000";
    tmp(76453) := x"0000";
    tmp(76454) := x"0000";
    tmp(76455) := x"0000";
    tmp(76456) := x"0000";
    tmp(76457) := x"0000";
    tmp(76458) := x"0000";
    tmp(76459) := x"0000";
    tmp(76460) := x"0000";
    tmp(76461) := x"0000";
    tmp(76462) := x"0000";
    tmp(76463) := x"0000";
    tmp(76464) := x"0000";
    tmp(76465) := x"0000";
    tmp(76466) := x"0000";
    tmp(76467) := x"0000";
    tmp(76468) := x"0000";
    tmp(76469) := x"0000";
    tmp(76470) := x"0000";
    tmp(76471) := x"0000";
    tmp(76472) := x"0000";
    tmp(76473) := x"0000";
    tmp(76474) := x"0000";
    tmp(76475) := x"0000";
    tmp(76476) := x"0000";
    tmp(76477) := x"0000";
    tmp(76478) := x"0000";
    tmp(76479) := x"0000";
    tmp(76480) := x"0000";
    tmp(76481) := x"0000";
    tmp(76482) := x"0000";
    tmp(76483) := x"0000";
    tmp(76484) := x"0000";
    tmp(76485) := x"0000";
    tmp(76486) := x"0000";
    tmp(76487) := x"0000";
    tmp(76488) := x"0000";
    tmp(76489) := x"0000";
    tmp(76490) := x"0000";
    tmp(76491) := x"0000";
    tmp(76492) := x"0000";
    tmp(76493) := x"0000";
    tmp(76494) := x"0000";
    tmp(76495) := x"0000";
    tmp(76496) := x"0000";
    tmp(76497) := x"0000";
    tmp(76498) := x"0000";
    tmp(76499) := x"0000";
    tmp(76500) := x"0000";
    tmp(76501) := x"0000";
    tmp(76502) := x"0000";
    tmp(76503) := x"0000";
    tmp(76504) := x"0000";
    tmp(76505) := x"0000";
    tmp(76506) := x"0000";
    tmp(76507) := x"0000";
    tmp(76508) := x"0000";
    tmp(76509) := x"0000";
    tmp(76510) := x"0000";
    tmp(76511) := x"0000";
    tmp(76512) := x"0000";
    tmp(76513) := x"0000";
    tmp(76514) := x"0000";
    tmp(76515) := x"0000";
    tmp(76516) := x"0000";
    tmp(76517) := x"0000";
    tmp(76518) := x"0000";
    tmp(76519) := x"0000";
    tmp(76520) := x"0000";
    tmp(76521) := x"0000";
    tmp(76522) := x"0000";
    tmp(76523) := x"0000";
    tmp(76524) := x"0000";
    tmp(76525) := x"0000";
    tmp(76526) := x"0000";
    tmp(76527) := x"0000";
    tmp(76528) := x"0000";
    tmp(76529) := x"0000";
    tmp(76530) := x"0000";
    tmp(76531) := x"0000";
    tmp(76532) := x"0000";
    tmp(76533) := x"0000";
    tmp(76534) := x"0000";
    tmp(76535) := x"0000";
    tmp(76536) := x"0000";
    tmp(76537) := x"0000";
    tmp(76538) := x"0000";
    tmp(76539) := x"0000";
    tmp(76540) := x"0000";
    tmp(76541) := x"0000";
    tmp(76542) := x"0000";
    tmp(76543) := x"0000";
    tmp(76544) := x"0000";
    tmp(76545) := x"0000";
    tmp(76546) := x"0000";
    tmp(76547) := x"0000";
    tmp(76548) := x"0000";
    tmp(76549) := x"0000";
    tmp(76550) := x"0000";
    tmp(76551) := x"0000";
    tmp(76552) := x"0000";
    tmp(76553) := x"0000";
    tmp(76554) := x"0000";
    tmp(76555) := x"0000";
    tmp(76556) := x"0000";
    tmp(76557) := x"0000";
    tmp(76558) := x"0000";
    tmp(76559) := x"0000";
    tmp(76560) := x"0000";
    tmp(76561) := x"0000";
    tmp(76562) := x"0000";
    tmp(76563) := x"0020";
    tmp(76564) := x"0020";
    tmp(76565) := x"0020";
    tmp(76566) := x"0040";
    tmp(76567) := x"0041";
    tmp(76568) := x"0041";
    tmp(76569) := x"0040";
    tmp(76570) := x"0040";
    tmp(76571) := x"0040";
    tmp(76572) := x"0040";
    tmp(76573) := x"0040";
    tmp(76574) := x"0040";
    tmp(76575) := x"0040";
    tmp(76576) := x"0040";
    tmp(76577) := x"0040";
    tmp(76578) := x"0040";
    tmp(76579) := x"0040";
    tmp(76580) := x"0040";
    tmp(76581) := x"0040";
    tmp(76582) := x"0040";
    tmp(76583) := x"0040";
    tmp(76584) := x"0040";
    tmp(76585) := x"0020";
    tmp(76586) := x"0020";
    tmp(76587) := x"0020";
    tmp(76588) := x"0020";
    tmp(76589) := x"0020";
    tmp(76590) := x"0020";
    tmp(76591) := x"0020";
    tmp(76592) := x"0020";
    tmp(76593) := x"0020";
    tmp(76594) := x"0020";
    tmp(76595) := x"0040";
    tmp(76596) := x"0040";
    tmp(76597) := x"0040";
    tmp(76598) := x"0040";
    tmp(76599) := x"0040";
    tmp(76600) := x"0020";
    tmp(76601) := x"0020";
    tmp(76602) := x"0020";
    tmp(76603) := x"0020";
    tmp(76604) := x"0020";
    tmp(76605) := x"0020";
    tmp(76606) := x"0820";
    tmp(76607) := x"0840";
    tmp(76608) := x"0040";
    tmp(76609) := x"0040";
    tmp(76610) := x"0040";
    tmp(76611) := x"0040";
    tmp(76612) := x"0040";
    tmp(76613) := x"0020";
    tmp(76614) := x"0020";
    tmp(76615) := x"0040";
    tmp(76616) := x"0040";
    tmp(76617) := x"0040";
    tmp(76618) := x"0820";
    tmp(76619) := x"0820";
    tmp(76620) := x"0820";
    tmp(76621) := x"1020";
    tmp(76622) := x"1020";
    tmp(76623) := x"1020";
    tmp(76624) := x"1020";
    tmp(76625) := x"1020";
    tmp(76626) := x"1020";
    tmp(76627) := x"1000";
    tmp(76628) := x"1000";
    tmp(76629) := x"1000";
    tmp(76630) := x"1000";
    tmp(76631) := x"1000";
    tmp(76632) := x"1000";
    tmp(76633) := x"1000";
    tmp(76634) := x"1000";
    tmp(76635) := x"1000";
    tmp(76636) := x"1000";
    tmp(76637) := x"1800";
    tmp(76638) := x"1000";
    tmp(76639) := x"1800";
    tmp(76640) := x"1800";
    tmp(76641) := x"1800";
    tmp(76642) := x"1800";
    tmp(76643) := x"2000";
    tmp(76644) := x"2020";
    tmp(76645) := x"2820";
    tmp(76646) := x"2020";
    tmp(76647) := x"2000";
    tmp(76648) := x"2020";
    tmp(76649) := x"2020";
    tmp(76650) := x"2000";
    tmp(76651) := x"1800";
    tmp(76652) := x"2020";
    tmp(76653) := x"2820";
    tmp(76654) := x"2020";
    tmp(76655) := x"2000";
    tmp(76656) := x"2000";
    tmp(76657) := x"2020";
    tmp(76658) := x"2020";
    tmp(76659) := x"2020";
    tmp(76660) := x"1800";
    tmp(76661) := x"1000";
    tmp(76662) := x"1000";
    tmp(76663) := x"1000";
    tmp(76664) := x"0800";
    tmp(76665) := x"0800";
    tmp(76666) := x"1000";
    tmp(76667) := x"1000";
    tmp(76668) := x"0820";
    tmp(76669) := x"0020";
    tmp(76670) := x"0020";
    tmp(76671) := x"0020";
    tmp(76672) := x"0020";
    tmp(76673) := x"0020";
    tmp(76674) := x"0020";
    tmp(76675) := x"0020";
    tmp(76676) := x"0000";
    tmp(76677) := x"0000";
    tmp(76678) := x"0000";
    tmp(76679) := x"0000";
    tmp(76680) := x"0000";
    tmp(76681) := x"0000";
    tmp(76682) := x"0000";
    tmp(76683) := x"0000";
    tmp(76684) := x"0000";
    tmp(76685) := x"0000";
    tmp(76686) := x"0000";
    tmp(76687) := x"0000";
    tmp(76688) := x"0000";
    tmp(76689) := x"0000";
    tmp(76690) := x"0000";
    tmp(76691) := x"0000";
    tmp(76692) := x"0000";
    tmp(76693) := x"0000";
    tmp(76694) := x"0000";
    tmp(76695) := x"0000";
    tmp(76696) := x"0000";
    tmp(76697) := x"0000";
    tmp(76698) := x"0000";
    tmp(76699) := x"0000";
    tmp(76700) := x"0000";
    tmp(76701) := x"0000";
    tmp(76702) := x"0000";
    tmp(76703) := x"0000";
    tmp(76704) := x"0000";
    tmp(76705) := x"0000";
    tmp(76706) := x"0000";
    tmp(76707) := x"0000";
    tmp(76708) := x"0000";
    tmp(76709) := x"0000";
    tmp(76710) := x"0000";
    tmp(76711) := x"0000";
    tmp(76712) := x"0000";
    tmp(76713) := x"0000";
    tmp(76714) := x"0000";
    tmp(76715) := x"0000";
    tmp(76716) := x"0000";
    tmp(76717) := x"0000";
    tmp(76718) := x"0000";
    tmp(76719) := x"0000";
    tmp(76720) := x"0000";
    tmp(76721) := x"0000";
    tmp(76722) := x"0000";
    tmp(76723) := x"0000";
    tmp(76724) := x"0000";
    tmp(76725) := x"0000";
    tmp(76726) := x"0000";
    tmp(76727) := x"0000";
    tmp(76728) := x"0000";
    tmp(76729) := x"0000";
    tmp(76730) := x"0000";
    tmp(76731) := x"0000";
    tmp(76732) := x"0000";
    tmp(76733) := x"0000";
    tmp(76734) := x"0000";
    tmp(76735) := x"0000";
    tmp(76736) := x"0000";
    tmp(76737) := x"0000";
    tmp(76738) := x"0000";
    tmp(76739) := x"0000";
    tmp(76740) := x"0000";
    tmp(76741) := x"0000";
    tmp(76742) := x"0000";
    tmp(76743) := x"0000";
    tmp(76744) := x"0000";
    tmp(76745) := x"0000";
    tmp(76746) := x"0000";
    tmp(76747) := x"0000";
    tmp(76748) := x"0000";
    tmp(76749) := x"0000";
    tmp(76750) := x"0000";
    tmp(76751) := x"0000";
    tmp(76752) := x"0000";
    tmp(76753) := x"0000";
    tmp(76754) := x"0000";
    tmp(76755) := x"0000";
    tmp(76756) := x"0000";
    tmp(76757) := x"0000";
    tmp(76758) := x"0000";
    tmp(76759) := x"0000";
    tmp(76760) := x"0000";
    tmp(76761) := x"0000";
    tmp(76762) := x"0000";
    tmp(76763) := x"0000";
    tmp(76764) := x"0000";
    tmp(76765) := x"0000";
    tmp(76766) := x"0000";
    tmp(76767) := x"0000";
    tmp(76768) := x"0000";
    tmp(76769) := x"0000";
    tmp(76770) := x"0000";
    tmp(76771) := x"0000";
    tmp(76772) := x"0000";
    tmp(76773) := x"0000";
    tmp(76774) := x"0000";
    tmp(76775) := x"0000";
    tmp(76776) := x"0000";
    tmp(76777) := x"0000";
    tmp(76778) := x"0000";
    tmp(76779) := x"0000";
    tmp(76780) := x"0000";
    tmp(76781) := x"0000";
    tmp(76782) := x"0000";
    tmp(76783) := x"0000";
    tmp(76784) := x"0000";
    tmp(76785) := x"0000";
    tmp(76786) := x"0000";
    tmp(76787) := x"0000";
    tmp(76788) := x"0000";
    tmp(76789) := x"0000";
    tmp(76790) := x"0000";
    tmp(76791) := x"0000";
    tmp(76792) := x"0000";
    tmp(76793) := x"0000";
    tmp(76794) := x"0000";
    tmp(76795) := x"0000";
    tmp(76796) := x"0000";
    tmp(76797) := x"0000";
    tmp(76798) := x"0000";
    tmp(76799) := x"0000";
    tmp(76800) := x"0000";
    tmp(76801) := x"0000";
    tmp(76802) := x"0000";
    tmp(76803) := x"0020";
    tmp(76804) := x"0020";
    tmp(76805) := x"0020";
    tmp(76806) := x"0020";
    tmp(76807) := x"0020";
    tmp(76808) := x"0041";
    tmp(76809) := x"0041";
    tmp(76810) := x"0040";
    tmp(76811) := x"0040";
    tmp(76812) := x"0040";
    tmp(76813) := x"0040";
    tmp(76814) := x"0040";
    tmp(76815) := x"0040";
    tmp(76816) := x"0040";
    tmp(76817) := x"0040";
    tmp(76818) := x"0040";
    tmp(76819) := x"0040";
    tmp(76820) := x"0040";
    tmp(76821) := x"0040";
    tmp(76822) := x"0040";
    tmp(76823) := x"0040";
    tmp(76824) := x"0040";
    tmp(76825) := x"0040";
    tmp(76826) := x"0020";
    tmp(76827) := x"0020";
    tmp(76828) := x"0020";
    tmp(76829) := x"0020";
    tmp(76830) := x"0020";
    tmp(76831) := x"0020";
    tmp(76832) := x"0020";
    tmp(76833) := x"0020";
    tmp(76834) := x"0020";
    tmp(76835) := x"0020";
    tmp(76836) := x"0020";
    tmp(76837) := x"0020";
    tmp(76838) := x"0040";
    tmp(76839) := x"0840";
    tmp(76840) := x"0840";
    tmp(76841) := x"0040";
    tmp(76842) := x"0040";
    tmp(76843) := x"0040";
    tmp(76844) := x"0020";
    tmp(76845) := x"0020";
    tmp(76846) := x"0020";
    tmp(76847) := x"0820";
    tmp(76848) := x"0820";
    tmp(76849) := x"0820";
    tmp(76850) := x"0820";
    tmp(76851) := x"0020";
    tmp(76852) := x"0040";
    tmp(76853) := x"0020";
    tmp(76854) := x"0020";
    tmp(76855) := x"0040";
    tmp(76856) := x"0040";
    tmp(76857) := x"0040";
    tmp(76858) := x"0020";
    tmp(76859) := x"0820";
    tmp(76860) := x"1020";
    tmp(76861) := x"1020";
    tmp(76862) := x"1020";
    tmp(76863) := x"1000";
    tmp(76864) := x"1800";
    tmp(76865) := x"1800";
    tmp(76866) := x"1800";
    tmp(76867) := x"1800";
    tmp(76868) := x"1800";
    tmp(76869) := x"1800";
    tmp(76870) := x"1800";
    tmp(76871) := x"1000";
    tmp(76872) := x"1000";
    tmp(76873) := x"0800";
    tmp(76874) := x"1000";
    tmp(76875) := x"1000";
    tmp(76876) := x"1800";
    tmp(76877) := x"1800";
    tmp(76878) := x"1800";
    tmp(76879) := x"1800";
    tmp(76880) := x"1800";
    tmp(76881) := x"1800";
    tmp(76882) := x"2000";
    tmp(76883) := x"2000";
    tmp(76884) := x"2820";
    tmp(76885) := x"2820";
    tmp(76886) := x"2020";
    tmp(76887) := x"2020";
    tmp(76888) := x"2020";
    tmp(76889) := x"2020";
    tmp(76890) := x"1800";
    tmp(76891) := x"1800";
    tmp(76892) := x"1800";
    tmp(76893) := x"2000";
    tmp(76894) := x"2020";
    tmp(76895) := x"2020";
    tmp(76896) := x"2020";
    tmp(76897) := x"1800";
    tmp(76898) := x"1800";
    tmp(76899) := x"1800";
    tmp(76900) := x"1820";
    tmp(76901) := x"1820";
    tmp(76902) := x"0800";
    tmp(76903) := x"0800";
    tmp(76904) := x"0800";
    tmp(76905) := x"1000";
    tmp(76906) := x"1000";
    tmp(76907) := x"1000";
    tmp(76908) := x"0820";
    tmp(76909) := x"0020";
    tmp(76910) := x"0020";
    tmp(76911) := x"0020";
    tmp(76912) := x"0020";
    tmp(76913) := x"0020";
    tmp(76914) := x"0020";
    tmp(76915) := x"0020";
    tmp(76916) := x"0000";
    tmp(76917) := x"0000";
    tmp(76918) := x"0000";
    tmp(76919) := x"0000";
    tmp(76920) := x"0000";
    tmp(76921) := x"0000";
    tmp(76922) := x"0000";
    tmp(76923) := x"0000";
    tmp(76924) := x"0000";
    tmp(76925) := x"0000";
    tmp(76926) := x"0000";
    tmp(76927) := x"0000";
    tmp(76928) := x"0000";
    tmp(76929) := x"0000";
    tmp(76930) := x"0000";
    tmp(76931) := x"0000";
    tmp(76932) := x"0000";
    tmp(76933) := x"0000";
    tmp(76934) := x"0000";
    tmp(76935) := x"0000";
    tmp(76936) := x"0000";
    tmp(76937) := x"0000";
    tmp(76938) := x"0000";
    tmp(76939) := x"0000";
    tmp(76940) := x"0000";
    tmp(76941) := x"0000";
    tmp(76942) := x"0000";
    tmp(76943) := x"0000";
    tmp(76944) := x"0000";
    tmp(76945) := x"0000";
    tmp(76946) := x"0000";
    tmp(76947) := x"0000";
    tmp(76948) := x"0000";
    tmp(76949) := x"0000";
    tmp(76950) := x"0000";
    tmp(76951) := x"0000";
    tmp(76952) := x"0000";
    tmp(76953) := x"0000";
    tmp(76954) := x"0000";
    tmp(76955) := x"0000";
    tmp(76956) := x"0000";
    tmp(76957) := x"0000";
    tmp(76958) := x"0000";
    tmp(76959) := x"0000";
    tmp(76960) := x"0000";
    tmp(76961) := x"0000";
    tmp(76962) := x"0000";
    tmp(76963) := x"0000";
    tmp(76964) := x"0000";
    tmp(76965) := x"0000";
    tmp(76966) := x"0000";
    tmp(76967) := x"0000";
    tmp(76968) := x"0000";
    tmp(76969) := x"0000";
    tmp(76970) := x"0000";
    tmp(76971) := x"0000";
    tmp(76972) := x"0000";
    tmp(76973) := x"0000";
    tmp(76974) := x"0000";
    tmp(76975) := x"0000";
    tmp(76976) := x"0000";
    tmp(76977) := x"0000";
    tmp(76978) := x"0000";
    tmp(76979) := x"0000";
    tmp(76980) := x"0000";
    tmp(76981) := x"0000";
    tmp(76982) := x"0000";
    tmp(76983) := x"0000";
    tmp(76984) := x"0000";
    tmp(76985) := x"0000";
    tmp(76986) := x"0000";
    tmp(76987) := x"0000";
    tmp(76988) := x"0000";
    tmp(76989) := x"0000";
    tmp(76990) := x"0000";
    tmp(76991) := x"0000";
    tmp(76992) := x"0000";
    tmp(76993) := x"0000";
    tmp(76994) := x"0000";
    tmp(76995) := x"0000";
    tmp(76996) := x"0000";
    tmp(76997) := x"0000";
    tmp(76998) := x"0000";
    tmp(76999) := x"0000";
    tmp(77000) := x"0000";
    tmp(77001) := x"0000";
    tmp(77002) := x"0000";
    tmp(77003) := x"0000";
    tmp(77004) := x"0000";
    tmp(77005) := x"0000";
    tmp(77006) := x"0000";
    tmp(77007) := x"0000";
    tmp(77008) := x"0000";
    tmp(77009) := x"0000";
    tmp(77010) := x"0000";
    tmp(77011) := x"0000";
    tmp(77012) := x"0000";
    tmp(77013) := x"0000";
    tmp(77014) := x"0000";
    tmp(77015) := x"0000";
    tmp(77016) := x"0000";
    tmp(77017) := x"0000";
    tmp(77018) := x"0000";
    tmp(77019) := x"0000";
    tmp(77020) := x"0000";
    tmp(77021) := x"0000";
    tmp(77022) := x"0000";
    tmp(77023) := x"0000";
    tmp(77024) := x"0000";
    tmp(77025) := x"0000";
    tmp(77026) := x"0000";
    tmp(77027) := x"0000";
    tmp(77028) := x"0000";
    tmp(77029) := x"0000";
    tmp(77030) := x"0000";
    tmp(77031) := x"0000";
    tmp(77032) := x"0000";
    tmp(77033) := x"0000";
    tmp(77034) := x"0000";
    tmp(77035) := x"0000";
    tmp(77036) := x"0000";
    tmp(77037) := x"0000";
    tmp(77038) := x"0000";
    tmp(77039) := x"0000";
    tmp(77040) := x"0000";
    tmp(77041) := x"0000";
    tmp(77042) := x"0000";
    tmp(77043) := x"0020";
    tmp(77044) := x"0020";
    tmp(77045) := x"0020";
    tmp(77046) := x"0020";
    tmp(77047) := x"0020";
    tmp(77048) := x"0020";
    tmp(77049) := x"0040";
    tmp(77050) := x"0040";
    tmp(77051) := x"0040";
    tmp(77052) := x"0040";
    tmp(77053) := x"0020";
    tmp(77054) := x"0020";
    tmp(77055) := x"0020";
    tmp(77056) := x"0020";
    tmp(77057) := x"0020";
    tmp(77058) := x"0020";
    tmp(77059) := x"0020";
    tmp(77060) := x"0020";
    tmp(77061) := x"0020";
    tmp(77062) := x"0020";
    tmp(77063) := x"0020";
    tmp(77064) := x"0020";
    tmp(77065) := x"0020";
    tmp(77066) := x"0020";
    tmp(77067) := x"0020";
    tmp(77068) := x"0020";
    tmp(77069) := x"0020";
    tmp(77070) := x"0020";
    tmp(77071) := x"0020";
    tmp(77072) := x"0020";
    tmp(77073) := x"0020";
    tmp(77074) := x"0020";
    tmp(77075) := x"0020";
    tmp(77076) := x"0020";
    tmp(77077) := x"0020";
    tmp(77078) := x"0020";
    tmp(77079) := x"0020";
    tmp(77080) := x"0020";
    tmp(77081) := x"0040";
    tmp(77082) := x"0040";
    tmp(77083) := x"0040";
    tmp(77084) := x"0020";
    tmp(77085) := x"0020";
    tmp(77086) := x"0020";
    tmp(77087) := x"0000";
    tmp(77088) := x"0800";
    tmp(77089) := x"0800";
    tmp(77090) := x"0820";
    tmp(77091) := x"0820";
    tmp(77092) := x"0820";
    tmp(77093) := x"0020";
    tmp(77094) := x"0020";
    tmp(77095) := x"0040";
    tmp(77096) := x"0040";
    tmp(77097) := x"0040";
    tmp(77098) := x"0020";
    tmp(77099) := x"0820";
    tmp(77100) := x"0820";
    tmp(77101) := x"1000";
    tmp(77102) := x"1000";
    tmp(77103) := x"1000";
    tmp(77104) := x"1800";
    tmp(77105) := x"1800";
    tmp(77106) := x"1800";
    tmp(77107) := x"1800";
    tmp(77108) := x"1800";
    tmp(77109) := x"1800";
    tmp(77110) := x"1800";
    tmp(77111) := x"1000";
    tmp(77112) := x"0800";
    tmp(77113) := x"0800";
    tmp(77114) := x"1000";
    tmp(77115) := x"1000";
    tmp(77116) := x"1000";
    tmp(77117) := x"1000";
    tmp(77118) := x"1800";
    tmp(77119) := x"1800";
    tmp(77120) := x"1800";
    tmp(77121) := x"1800";
    tmp(77122) := x"1800";
    tmp(77123) := x"2000";
    tmp(77124) := x"2020";
    tmp(77125) := x"2820";
    tmp(77126) := x"2820";
    tmp(77127) := x"2820";
    tmp(77128) := x"2020";
    tmp(77129) := x"1000";
    tmp(77130) := x"1000";
    tmp(77131) := x"2020";
    tmp(77132) := x"2820";
    tmp(77133) := x"2020";
    tmp(77134) := x"1820";
    tmp(77135) := x"1000";
    tmp(77136) := x"1000";
    tmp(77137) := x"1820";
    tmp(77138) := x"1820";
    tmp(77139) := x"1000";
    tmp(77140) := x"0800";
    tmp(77141) := x"0800";
    tmp(77142) := x"0800";
    tmp(77143) := x"0800";
    tmp(77144) := x"0800";
    tmp(77145) := x"1000";
    tmp(77146) := x"1000";
    tmp(77147) := x"0820";
    tmp(77148) := x"0020";
    tmp(77149) := x"0020";
    tmp(77150) := x"0020";
    tmp(77151) := x"0020";
    tmp(77152) := x"0020";
    tmp(77153) := x"0020";
    tmp(77154) := x"0020";
    tmp(77155) := x"0020";
    tmp(77156) := x"0000";
    tmp(77157) := x"0000";
    tmp(77158) := x"0000";
    tmp(77159) := x"0000";
    tmp(77160) := x"0000";
    tmp(77161) := x"0000";
    tmp(77162) := x"0000";
    tmp(77163) := x"0000";
    tmp(77164) := x"0000";
    tmp(77165) := x"0000";
    tmp(77166) := x"0000";
    tmp(77167) := x"0000";
    tmp(77168) := x"0000";
    tmp(77169) := x"0000";
    tmp(77170) := x"0000";
    tmp(77171) := x"0000";
    tmp(77172) := x"0000";
    tmp(77173) := x"0000";
    tmp(77174) := x"0000";
    tmp(77175) := x"0000";
    tmp(77176) := x"0000";
    tmp(77177) := x"0000";
    tmp(77178) := x"0000";
    tmp(77179) := x"0000";
    tmp(77180) := x"0000";
    tmp(77181) := x"0000";
    tmp(77182) := x"0000";
    tmp(77183) := x"0000";
    tmp(77184) := x"0000";
    tmp(77185) := x"0000";
    tmp(77186) := x"0000";
    tmp(77187) := x"0000";
    tmp(77188) := x"0000";
    tmp(77189) := x"0000";
    tmp(77190) := x"0000";
    tmp(77191) := x"0000";
    tmp(77192) := x"0000";
    tmp(77193) := x"0000";
    tmp(77194) := x"0000";
    tmp(77195) := x"0000";
    tmp(77196) := x"0000";
    tmp(77197) := x"0000";
    tmp(77198) := x"0000";
    tmp(77199) := x"0000";
    tmp(77200) := x"0000";
    tmp(77201) := x"0000";
    tmp(77202) := x"0000";
    tmp(77203) := x"0000";
    tmp(77204) := x"0000";
    tmp(77205) := x"0000";
    tmp(77206) := x"0000";
    tmp(77207) := x"0000";
    tmp(77208) := x"0000";
    tmp(77209) := x"0000";
    tmp(77210) := x"0000";
    tmp(77211) := x"0000";
    tmp(77212) := x"0000";
    tmp(77213) := x"0000";
    tmp(77214) := x"0000";
    tmp(77215) := x"0000";
    tmp(77216) := x"0000";
    tmp(77217) := x"0000";
    tmp(77218) := x"0000";
    tmp(77219) := x"0000";
    tmp(77220) := x"0000";
    tmp(77221) := x"0000";
    tmp(77222) := x"0000";
    tmp(77223) := x"0000";
    tmp(77224) := x"0000";
    tmp(77225) := x"0000";
    tmp(77226) := x"0000";
    tmp(77227) := x"0000";
    tmp(77228) := x"0000";
    tmp(77229) := x"0000";
    tmp(77230) := x"0000";
    tmp(77231) := x"0000";
    tmp(77232) := x"0000";
    tmp(77233) := x"0000";
    tmp(77234) := x"0000";
    tmp(77235) := x"0000";
    tmp(77236) := x"0000";
    tmp(77237) := x"0000";
    tmp(77238) := x"0000";
    tmp(77239) := x"0000";
    tmp(77240) := x"0000";
    tmp(77241) := x"0000";
    tmp(77242) := x"0000";
    tmp(77243) := x"0000";
    tmp(77244) := x"0000";
    tmp(77245) := x"0000";
    tmp(77246) := x"0000";
    tmp(77247) := x"0000";
    tmp(77248) := x"0000";
    tmp(77249) := x"0000";
    tmp(77250) := x"0000";
    tmp(77251) := x"0000";
    tmp(77252) := x"0000";
    tmp(77253) := x"0000";
    tmp(77254) := x"0000";
    tmp(77255) := x"0000";
    tmp(77256) := x"0000";
    tmp(77257) := x"0000";
    tmp(77258) := x"0000";
    tmp(77259) := x"0000";
    tmp(77260) := x"0000";
    tmp(77261) := x"0000";
    tmp(77262) := x"0000";
    tmp(77263) := x"0000";
    tmp(77264) := x"0000";
    tmp(77265) := x"0000";
    tmp(77266) := x"0000";
    tmp(77267) := x"0000";
    tmp(77268) := x"0000";
    tmp(77269) := x"0000";
    tmp(77270) := x"0000";
    tmp(77271) := x"0000";
    tmp(77272) := x"0000";
    tmp(77273) := x"0000";
    tmp(77274) := x"0000";
    tmp(77275) := x"0000";
    tmp(77276) := x"0000";
    tmp(77277) := x"0000";
    tmp(77278) := x"0000";
    tmp(77279) := x"0000";
    tmp(77280) := x"0000";
    tmp(77281) := x"0000";
    tmp(77282) := x"0000";
    tmp(77283) := x"0020";
    tmp(77284) := x"0020";
    tmp(77285) := x"0020";
    tmp(77286) := x"0020";
    tmp(77287) := x"0020";
    tmp(77288) := x"0020";
    tmp(77289) := x"0020";
    tmp(77290) := x"0020";
    tmp(77291) := x"0020";
    tmp(77292) := x"0020";
    tmp(77293) := x"0040";
    tmp(77294) := x"0040";
    tmp(77295) := x"0040";
    tmp(77296) := x"0020";
    tmp(77297) := x"0020";
    tmp(77298) := x"0040";
    tmp(77299) := x"0040";
    tmp(77300) := x"0040";
    tmp(77301) := x"0020";
    tmp(77302) := x"0020";
    tmp(77303) := x"0020";
    tmp(77304) := x"0020";
    tmp(77305) := x"0020";
    tmp(77306) := x"0020";
    tmp(77307) := x"0020";
    tmp(77308) := x"0020";
    tmp(77309) := x"0020";
    tmp(77310) := x"0020";
    tmp(77311) := x"0020";
    tmp(77312) := x"0020";
    tmp(77313) := x"0020";
    tmp(77314) := x"0020";
    tmp(77315) := x"0000";
    tmp(77316) := x"0000";
    tmp(77317) := x"0000";
    tmp(77318) := x"0000";
    tmp(77319) := x"0000";
    tmp(77320) := x"0000";
    tmp(77321) := x"0000";
    tmp(77322) := x"0020";
    tmp(77323) := x"0040";
    tmp(77324) := x"0040";
    tmp(77325) := x"0040";
    tmp(77326) := x"0020";
    tmp(77327) := x"0020";
    tmp(77328) := x"0000";
    tmp(77329) := x"0000";
    tmp(77330) := x"0800";
    tmp(77331) := x"0800";
    tmp(77332) := x"0820";
    tmp(77333) := x"0820";
    tmp(77334) := x"0820";
    tmp(77335) := x"0020";
    tmp(77336) := x"0020";
    tmp(77337) := x"0020";
    tmp(77338) := x"0020";
    tmp(77339) := x"0820";
    tmp(77340) := x"0800";
    tmp(77341) := x"0800";
    tmp(77342) := x"1000";
    tmp(77343) := x"1000";
    tmp(77344) := x"1000";
    tmp(77345) := x"1000";
    tmp(77346) := x"1000";
    tmp(77347) := x"1800";
    tmp(77348) := x"1800";
    tmp(77349) := x"1800";
    tmp(77350) := x"1800";
    tmp(77351) := x"1000";
    tmp(77352) := x"0800";
    tmp(77353) := x"0800";
    tmp(77354) := x"1000";
    tmp(77355) := x"1000";
    tmp(77356) := x"1000";
    tmp(77357) := x"1000";
    tmp(77358) := x"1800";
    tmp(77359) := x"1800";
    tmp(77360) := x"1820";
    tmp(77361) := x"1820";
    tmp(77362) := x"1820";
    tmp(77363) := x"1800";
    tmp(77364) := x"2020";
    tmp(77365) := x"2820";
    tmp(77366) := x"2820";
    tmp(77367) := x"2020";
    tmp(77368) := x"1800";
    tmp(77369) := x"1800";
    tmp(77370) := x"2020";
    tmp(77371) := x"2820";
    tmp(77372) := x"1820";
    tmp(77373) := x"0800";
    tmp(77374) := x"0800";
    tmp(77375) := x"1000";
    tmp(77376) := x"1000";
    tmp(77377) := x"0800";
    tmp(77378) := x"0800";
    tmp(77379) := x"0800";
    tmp(77380) := x"0800";
    tmp(77381) := x"0800";
    tmp(77382) := x"1000";
    tmp(77383) := x"0800";
    tmp(77384) := x"1000";
    tmp(77385) := x"1000";
    tmp(77386) := x"1000";
    tmp(77387) := x"0820";
    tmp(77388) := x"0020";
    tmp(77389) := x"0020";
    tmp(77390) := x"0020";
    tmp(77391) := x"0020";
    tmp(77392) := x"0020";
    tmp(77393) := x"0020";
    tmp(77394) := x"0020";
    tmp(77395) := x"0020";
    tmp(77396) := x"0020";
    tmp(77397) := x"0000";
    tmp(77398) := x"0000";
    tmp(77399) := x"0000";
    tmp(77400) := x"0000";
    tmp(77401) := x"0000";
    tmp(77402) := x"0000";
    tmp(77403) := x"0000";
    tmp(77404) := x"0000";
    tmp(77405) := x"0000";
    tmp(77406) := x"0000";
    tmp(77407) := x"0000";
    tmp(77408) := x"0000";
    tmp(77409) := x"0000";
    tmp(77410) := x"0000";
    tmp(77411) := x"0000";
    tmp(77412) := x"0000";
    tmp(77413) := x"0000";
    tmp(77414) := x"0000";
    tmp(77415) := x"0000";
    tmp(77416) := x"0000";
    tmp(77417) := x"0000";
    tmp(77418) := x"0000";
    tmp(77419) := x"0000";
    tmp(77420) := x"0000";
    tmp(77421) := x"0000";
    tmp(77422) := x"0000";
    tmp(77423) := x"0000";
    tmp(77424) := x"0000";
    tmp(77425) := x"0000";
    tmp(77426) := x"0000";
    tmp(77427) := x"0000";
    tmp(77428) := x"0000";
    tmp(77429) := x"0000";
    tmp(77430) := x"0000";
    tmp(77431) := x"0000";
    tmp(77432) := x"0000";
    tmp(77433) := x"0000";
    tmp(77434) := x"0000";
    tmp(77435) := x"0000";
    tmp(77436) := x"0000";
    tmp(77437) := x"0000";
    tmp(77438) := x"0000";
    tmp(77439) := x"0000";
    tmp(77440) := x"0000";
    tmp(77441) := x"0000";
    tmp(77442) := x"0000";
    tmp(77443) := x"0000";
    tmp(77444) := x"0000";
    tmp(77445) := x"0000";
    tmp(77446) := x"0000";
    tmp(77447) := x"0000";
    tmp(77448) := x"0000";
    tmp(77449) := x"0000";
    tmp(77450) := x"0000";
    tmp(77451) := x"0000";
    tmp(77452) := x"0000";
    tmp(77453) := x"0000";
    tmp(77454) := x"0000";
    tmp(77455) := x"0000";
    tmp(77456) := x"0000";
    tmp(77457) := x"0000";
    tmp(77458) := x"0000";
    tmp(77459) := x"0000";
    tmp(77460) := x"0000";
    tmp(77461) := x"0000";
    tmp(77462) := x"0000";
    tmp(77463) := x"0000";
    tmp(77464) := x"0000";
    tmp(77465) := x"0000";
    tmp(77466) := x"0000";
    tmp(77467) := x"0000";
    tmp(77468) := x"0000";
    tmp(77469) := x"0000";
    tmp(77470) := x"0000";
    tmp(77471) := x"0000";
    tmp(77472) := x"0000";
    tmp(77473) := x"0000";
    tmp(77474) := x"0000";
    tmp(77475) := x"0000";
    tmp(77476) := x"0000";
    tmp(77477) := x"0000";
    tmp(77478) := x"0000";
    tmp(77479) := x"0000";
    tmp(77480) := x"0000";
    tmp(77481) := x"0000";
    tmp(77482) := x"0000";
    tmp(77483) := x"0000";
    tmp(77484) := x"0000";
    tmp(77485) := x"0000";
    tmp(77486) := x"0000";
    tmp(77487) := x"0000";
    tmp(77488) := x"0000";
    tmp(77489) := x"0000";
    tmp(77490) := x"0000";
    tmp(77491) := x"0000";
    tmp(77492) := x"0000";
    tmp(77493) := x"0000";
    tmp(77494) := x"0000";
    tmp(77495) := x"0000";
    tmp(77496) := x"0000";
    tmp(77497) := x"0000";
    tmp(77498) := x"0000";
    tmp(77499) := x"0000";
    tmp(77500) := x"0000";
    tmp(77501) := x"0000";
    tmp(77502) := x"0000";
    tmp(77503) := x"0000";
    tmp(77504) := x"0000";
    tmp(77505) := x"0000";
    tmp(77506) := x"0000";
    tmp(77507) := x"0000";
    tmp(77508) := x"0000";
    tmp(77509) := x"0000";
    tmp(77510) := x"0000";
    tmp(77511) := x"0000";
    tmp(77512) := x"0000";
    tmp(77513) := x"0000";
    tmp(77514) := x"0000";
    tmp(77515) := x"0000";
    tmp(77516) := x"0000";
    tmp(77517) := x"0000";
    tmp(77518) := x"0000";
    tmp(77519) := x"0000";
    tmp(77520) := x"0000";
    tmp(77521) := x"0000";
    tmp(77522) := x"0000";
    tmp(77523) := x"0000";
    tmp(77524) := x"0020";
    tmp(77525) := x"0020";
    tmp(77526) := x"0020";
    tmp(77527) := x"0020";
    tmp(77528) := x"0020";
    tmp(77529) := x"0020";
    tmp(77530) := x"0020";
    tmp(77531) := x"0020";
    tmp(77532) := x"0040";
    tmp(77533) := x"0041";
    tmp(77534) := x"0041";
    tmp(77535) := x"0040";
    tmp(77536) := x"0040";
    tmp(77537) := x"0040";
    tmp(77538) := x"0040";
    tmp(77539) := x"0040";
    tmp(77540) := x"0040";
    tmp(77541) := x"0040";
    tmp(77542) := x"0040";
    tmp(77543) := x"0040";
    tmp(77544) := x"0040";
    tmp(77545) := x"0040";
    tmp(77546) := x"0020";
    tmp(77547) := x"0020";
    tmp(77548) := x"0020";
    tmp(77549) := x"0040";
    tmp(77550) := x"0040";
    tmp(77551) := x"0020";
    tmp(77552) := x"0020";
    tmp(77553) := x"0020";
    tmp(77554) := x"0020";
    tmp(77555) := x"0020";
    tmp(77556) := x"0020";
    tmp(77557) := x"0020";
    tmp(77558) := x"0000";
    tmp(77559) := x"0000";
    tmp(77560) := x"0000";
    tmp(77561) := x"0000";
    tmp(77562) := x"0000";
    tmp(77563) := x"0000";
    tmp(77564) := x"0020";
    tmp(77565) := x"0020";
    tmp(77566) := x"0020";
    tmp(77567) := x"0020";
    tmp(77568) := x"0000";
    tmp(77569) := x"0000";
    tmp(77570) := x"0000";
    tmp(77571) := x"0800";
    tmp(77572) := x"0800";
    tmp(77573) := x"0800";
    tmp(77574) := x"0820";
    tmp(77575) := x"0820";
    tmp(77576) := x"0820";
    tmp(77577) := x"0020";
    tmp(77578) := x"0020";
    tmp(77579) := x"0820";
    tmp(77580) := x"0800";
    tmp(77581) := x"0800";
    tmp(77582) := x"0800";
    tmp(77583) := x"1000";
    tmp(77584) := x"1000";
    tmp(77585) := x"1000";
    tmp(77586) := x"1000";
    tmp(77587) := x"1800";
    tmp(77588) := x"1800";
    tmp(77589) := x"1800";
    tmp(77590) := x"1000";
    tmp(77591) := x"0800";
    tmp(77592) := x"0800";
    tmp(77593) := x"1000";
    tmp(77594) := x"1000";
    tmp(77595) := x"1000";
    tmp(77596) := x"1000";
    tmp(77597) := x"1000";
    tmp(77598) := x"1000";
    tmp(77599) := x"1800";
    tmp(77600) := x"1000";
    tmp(77601) := x"1000";
    tmp(77602) := x"1000";
    tmp(77603) := x"1000";
    tmp(77604) := x"2000";
    tmp(77605) := x"2820";
    tmp(77606) := x"2820";
    tmp(77607) := x"1800";
    tmp(77608) := x"1800";
    tmp(77609) := x"2820";
    tmp(77610) := x"2020";
    tmp(77611) := x"1000";
    tmp(77612) := x"0800";
    tmp(77613) := x"0800";
    tmp(77614) := x"1000";
    tmp(77615) := x"1000";
    tmp(77616) := x"1000";
    tmp(77617) := x"1020";
    tmp(77618) := x"0800";
    tmp(77619) := x"0000";
    tmp(77620) := x"0000";
    tmp(77621) := x"0800";
    tmp(77622) := x"1000";
    tmp(77623) := x"1000";
    tmp(77624) := x"0800";
    tmp(77625) := x"1000";
    tmp(77626) := x"0820";
    tmp(77627) := x"0020";
    tmp(77628) := x"0020";
    tmp(77629) := x"0020";
    tmp(77630) := x"0020";
    tmp(77631) := x"0020";
    tmp(77632) := x"0020";
    tmp(77633) := x"0020";
    tmp(77634) := x"0020";
    tmp(77635) := x"0020";
    tmp(77636) := x"0000";
    tmp(77637) := x"0000";
    tmp(77638) := x"0000";
    tmp(77639) := x"0000";
    tmp(77640) := x"0000";
    tmp(77641) := x"0000";
    tmp(77642) := x"0000";
    tmp(77643) := x"0000";
    tmp(77644) := x"0000";
    tmp(77645) := x"0000";
    tmp(77646) := x"0000";
    tmp(77647) := x"0000";
    tmp(77648) := x"0000";
    tmp(77649) := x"0000";
    tmp(77650) := x"0000";
    tmp(77651) := x"0000";
    tmp(77652) := x"0000";
    tmp(77653) := x"0000";
    tmp(77654) := x"0000";
    tmp(77655) := x"0000";
    tmp(77656) := x"0000";
    tmp(77657) := x"0000";
    tmp(77658) := x"0000";
    tmp(77659) := x"0000";
    tmp(77660) := x"0000";
    tmp(77661) := x"0000";
    tmp(77662) := x"0000";
    tmp(77663) := x"0000";
    tmp(77664) := x"0000";
    tmp(77665) := x"0000";
    tmp(77666) := x"0000";
    tmp(77667) := x"0000";
    tmp(77668) := x"0000";
    tmp(77669) := x"0000";
    tmp(77670) := x"0000";
    tmp(77671) := x"0000";
    tmp(77672) := x"0000";
    tmp(77673) := x"0000";
    tmp(77674) := x"0000";
    tmp(77675) := x"0000";
    tmp(77676) := x"0000";
    tmp(77677) := x"0000";
    tmp(77678) := x"0000";
    tmp(77679) := x"0000";
    tmp(77680) := x"0000";
    tmp(77681) := x"0000";
    tmp(77682) := x"0000";
    tmp(77683) := x"0000";
    tmp(77684) := x"0000";
    tmp(77685) := x"0000";
    tmp(77686) := x"0000";
    tmp(77687) := x"0000";
    tmp(77688) := x"0000";
    tmp(77689) := x"0000";
    tmp(77690) := x"0000";
    tmp(77691) := x"0000";
    tmp(77692) := x"0000";
    tmp(77693) := x"0000";
    tmp(77694) := x"0000";
    tmp(77695) := x"0000";
    tmp(77696) := x"0000";
    tmp(77697) := x"0000";
    tmp(77698) := x"0000";
    tmp(77699) := x"0000";
    tmp(77700) := x"0000";
    tmp(77701) := x"0000";
    tmp(77702) := x"0000";
    tmp(77703) := x"0000";
    tmp(77704) := x"0000";
    tmp(77705) := x"0000";
    tmp(77706) := x"0000";
    tmp(77707) := x"0000";
    tmp(77708) := x"0000";
    tmp(77709) := x"0000";
    tmp(77710) := x"0000";
    tmp(77711) := x"0000";
    tmp(77712) := x"0000";
    tmp(77713) := x"0000";
    tmp(77714) := x"0000";
    tmp(77715) := x"0000";
    tmp(77716) := x"0000";
    tmp(77717) := x"0000";
    tmp(77718) := x"0000";
    tmp(77719) := x"0000";
    tmp(77720) := x"0000";
    tmp(77721) := x"0000";
    tmp(77722) := x"0000";
    tmp(77723) := x"0000";
    tmp(77724) := x"0000";
    tmp(77725) := x"0000";
    tmp(77726) := x"0000";
    tmp(77727) := x"0000";
    tmp(77728) := x"0000";
    tmp(77729) := x"0000";
    tmp(77730) := x"0000";
    tmp(77731) := x"0000";
    tmp(77732) := x"0000";
    tmp(77733) := x"0000";
    tmp(77734) := x"0000";
    tmp(77735) := x"0000";
    tmp(77736) := x"0000";
    tmp(77737) := x"0000";
    tmp(77738) := x"0000";
    tmp(77739) := x"0000";
    tmp(77740) := x"0000";
    tmp(77741) := x"0000";
    tmp(77742) := x"0000";
    tmp(77743) := x"0000";
    tmp(77744) := x"0000";
    tmp(77745) := x"0000";
    tmp(77746) := x"0000";
    tmp(77747) := x"0000";
    tmp(77748) := x"0000";
    tmp(77749) := x"0000";
    tmp(77750) := x"0000";
    tmp(77751) := x"0000";
    tmp(77752) := x"0000";
    tmp(77753) := x"0000";
    tmp(77754) := x"0000";
    tmp(77755) := x"0000";
    tmp(77756) := x"0000";
    tmp(77757) := x"0000";
    tmp(77758) := x"0000";
    tmp(77759) := x"0000";
    tmp(77760) := x"0000";
    tmp(77761) := x"0000";
    tmp(77762) := x"0000";
    tmp(77763) := x"0000";
    tmp(77764) := x"0000";
    tmp(77765) := x"0020";
    tmp(77766) := x"0020";
    tmp(77767) := x"0020";
    tmp(77768) := x"0020";
    tmp(77769) := x"0020";
    tmp(77770) := x"0020";
    tmp(77771) := x"0020";
    tmp(77772) := x"0040";
    tmp(77773) := x"0040";
    tmp(77774) := x"0040";
    tmp(77775) := x"0040";
    tmp(77776) := x"0040";
    tmp(77777) := x"0040";
    tmp(77778) := x"0040";
    tmp(77779) := x"0040";
    tmp(77780) := x"0040";
    tmp(77781) := x"0040";
    tmp(77782) := x"0040";
    tmp(77783) := x"0040";
    tmp(77784) := x"0040";
    tmp(77785) := x"0040";
    tmp(77786) := x"0040";
    tmp(77787) := x"0040";
    tmp(77788) := x"0040";
    tmp(77789) := x"0040";
    tmp(77790) := x"0040";
    tmp(77791) := x"0040";
    tmp(77792) := x"0040";
    tmp(77793) := x"0040";
    tmp(77794) := x"0040";
    tmp(77795) := x"0040";
    tmp(77796) := x"0040";
    tmp(77797) := x"0040";
    tmp(77798) := x"0040";
    tmp(77799) := x"0040";
    tmp(77800) := x"0040";
    tmp(77801) := x"0040";
    tmp(77802) := x"0020";
    tmp(77803) := x"0020";
    tmp(77804) := x"0020";
    tmp(77805) := x"0021";
    tmp(77806) := x"0020";
    tmp(77807) := x"0020";
    tmp(77808) := x"0020";
    tmp(77809) := x"0000";
    tmp(77810) := x"0800";
    tmp(77811) := x"0800";
    tmp(77812) := x"0800";
    tmp(77813) := x"0800";
    tmp(77814) := x"1000";
    tmp(77815) := x"1020";
    tmp(77816) := x"0820";
    tmp(77817) := x"0820";
    tmp(77818) := x"0800";
    tmp(77819) := x"0800";
    tmp(77820) := x"0800";
    tmp(77821) := x"0800";
    tmp(77822) := x"0800";
    tmp(77823) := x"1000";
    tmp(77824) := x"1000";
    tmp(77825) := x"1000";
    tmp(77826) := x"1000";
    tmp(77827) := x"1000";
    tmp(77828) := x"1800";
    tmp(77829) := x"1000";
    tmp(77830) := x"1000";
    tmp(77831) := x"0800";
    tmp(77832) := x"1000";
    tmp(77833) := x"1000";
    tmp(77834) := x"1800";
    tmp(77835) := x"1800";
    tmp(77836) := x"1800";
    tmp(77837) := x"1000";
    tmp(77838) := x"1000";
    tmp(77839) := x"1000";
    tmp(77840) := x"1000";
    tmp(77841) := x"1000";
    tmp(77842) := x"1000";
    tmp(77843) := x"1800";
    tmp(77844) := x"2000";
    tmp(77845) := x"2820";
    tmp(77846) := x"2020";
    tmp(77847) := x"1000";
    tmp(77848) := x"1000";
    tmp(77849) := x"1000";
    tmp(77850) := x"0800";
    tmp(77851) := x"0800";
    tmp(77852) := x"0800";
    tmp(77853) := x"1000";
    tmp(77854) := x"1800";
    tmp(77855) := x"2020";
    tmp(77856) := x"0800";
    tmp(77857) := x"0000";
    tmp(77858) := x"0000";
    tmp(77859) := x"0800";
    tmp(77860) := x"0800";
    tmp(77861) := x"0800";
    tmp(77862) := x"1000";
    tmp(77863) := x"0800";
    tmp(77864) := x"0800";
    tmp(77865) := x"0820";
    tmp(77866) := x"0020";
    tmp(77867) := x"0020";
    tmp(77868) := x"0020";
    tmp(77869) := x"0020";
    tmp(77870) := x"0020";
    tmp(77871) := x"0020";
    tmp(77872) := x"0020";
    tmp(77873) := x"0020";
    tmp(77874) := x"0000";
    tmp(77875) := x"0000";
    tmp(77876) := x"0000";
    tmp(77877) := x"0000";
    tmp(77878) := x"0000";
    tmp(77879) := x"0000";
    tmp(77880) := x"0000";
    tmp(77881) := x"0000";
    tmp(77882) := x"0000";
    tmp(77883) := x"0000";
    tmp(77884) := x"0000";
    tmp(77885) := x"0000";
    tmp(77886) := x"0000";
    tmp(77887) := x"0000";
    tmp(77888) := x"0000";
    tmp(77889) := x"0000";
    tmp(77890) := x"0000";
    tmp(77891) := x"0000";
    tmp(77892) := x"0000";
    tmp(77893) := x"0000";
    tmp(77894) := x"0000";
    tmp(77895) := x"0000";
    tmp(77896) := x"0000";
    tmp(77897) := x"0000";
    tmp(77898) := x"0000";
    tmp(77899) := x"0000";
    tmp(77900) := x"0000";
    tmp(77901) := x"0000";
    tmp(77902) := x"0000";
    tmp(77903) := x"0000";
    tmp(77904) := x"0000";
    tmp(77905) := x"0000";
    tmp(77906) := x"0000";
    tmp(77907) := x"0000";
    tmp(77908) := x"0000";
    tmp(77909) := x"0000";
    tmp(77910) := x"0000";
    tmp(77911) := x"0000";
    tmp(77912) := x"0000";
    tmp(77913) := x"0000";
    tmp(77914) := x"0000";
    tmp(77915) := x"0000";
    tmp(77916) := x"0000";
    tmp(77917) := x"0000";
    tmp(77918) := x"0000";
    tmp(77919) := x"0000";
    tmp(77920) := x"0000";
    tmp(77921) := x"0000";
    tmp(77922) := x"0000";
    tmp(77923) := x"0000";
    tmp(77924) := x"0000";
    tmp(77925) := x"0000";
    tmp(77926) := x"0000";
    tmp(77927) := x"0000";
    tmp(77928) := x"0000";
    tmp(77929) := x"0000";
    tmp(77930) := x"0000";
    tmp(77931) := x"0000";
    tmp(77932) := x"0000";
    tmp(77933) := x"0000";
    tmp(77934) := x"0000";
    tmp(77935) := x"0000";
    tmp(77936) := x"0000";
    tmp(77937) := x"0000";
    tmp(77938) := x"0000";
    tmp(77939) := x"0000";
    tmp(77940) := x"0000";
    tmp(77941) := x"0000";
    tmp(77942) := x"0000";
    tmp(77943) := x"0000";
    tmp(77944) := x"0000";
    tmp(77945) := x"0000";
    tmp(77946) := x"0000";
    tmp(77947) := x"0000";
    tmp(77948) := x"0000";
    tmp(77949) := x"0000";
    tmp(77950) := x"0000";
    tmp(77951) := x"0000";
    tmp(77952) := x"0000";
    tmp(77953) := x"0000";
    tmp(77954) := x"0000";
    tmp(77955) := x"0000";
    tmp(77956) := x"0000";
    tmp(77957) := x"0000";
    tmp(77958) := x"0000";
    tmp(77959) := x"0000";
    tmp(77960) := x"0000";
    tmp(77961) := x"0000";
    tmp(77962) := x"0000";
    tmp(77963) := x"0000";
    tmp(77964) := x"0000";
    tmp(77965) := x"0000";
    tmp(77966) := x"0000";
    tmp(77967) := x"0000";
    tmp(77968) := x"0000";
    tmp(77969) := x"0000";
    tmp(77970) := x"0000";
    tmp(77971) := x"0000";
    tmp(77972) := x"0000";
    tmp(77973) := x"0000";
    tmp(77974) := x"0000";
    tmp(77975) := x"0000";
    tmp(77976) := x"0000";
    tmp(77977) := x"0000";
    tmp(77978) := x"0000";
    tmp(77979) := x"0000";
    tmp(77980) := x"0000";
    tmp(77981) := x"0000";
    tmp(77982) := x"0000";
    tmp(77983) := x"0000";
    tmp(77984) := x"0000";
    tmp(77985) := x"0000";
    tmp(77986) := x"0000";
    tmp(77987) := x"0000";
    tmp(77988) := x"0000";
    tmp(77989) := x"0000";
    tmp(77990) := x"0000";
    tmp(77991) := x"0000";
    tmp(77992) := x"0000";
    tmp(77993) := x"0000";
    tmp(77994) := x"0000";
    tmp(77995) := x"0000";
    tmp(77996) := x"0000";
    tmp(77997) := x"0000";
    tmp(77998) := x"0000";
    tmp(77999) := x"0000";
    tmp(78000) := x"0000";
    tmp(78001) := x"0000";
    tmp(78002) := x"0000";
    tmp(78003) := x"0000";
    tmp(78004) := x"0000";
    tmp(78005) := x"0000";
    tmp(78006) := x"0020";
    tmp(78007) := x"0020";
    tmp(78008) := x"0020";
    tmp(78009) := x"0020";
    tmp(78010) := x"0020";
    tmp(78011) := x"0020";
    tmp(78012) := x"0020";
    tmp(78013) := x"0040";
    tmp(78014) := x"0040";
    tmp(78015) := x"0040";
    tmp(78016) := x"0040";
    tmp(78017) := x"0040";
    tmp(78018) := x"0040";
    tmp(78019) := x"0040";
    tmp(78020) := x"0040";
    tmp(78021) := x"0040";
    tmp(78022) := x"0040";
    tmp(78023) := x"0040";
    tmp(78024) := x"0040";
    tmp(78025) := x"0040";
    tmp(78026) := x"0040";
    tmp(78027) := x"0040";
    tmp(78028) := x"0040";
    tmp(78029) := x"0040";
    tmp(78030) := x"0040";
    tmp(78031) := x"0040";
    tmp(78032) := x"0040";
    tmp(78033) := x"0040";
    tmp(78034) := x"0040";
    tmp(78035) := x"0040";
    tmp(78036) := x"0040";
    tmp(78037) := x"0040";
    tmp(78038) := x"0040";
    tmp(78039) := x"0040";
    tmp(78040) := x"0040";
    tmp(78041) := x"0041";
    tmp(78042) := x"0020";
    tmp(78043) := x"0021";
    tmp(78044) := x"0021";
    tmp(78045) := x"0021";
    tmp(78046) := x"0021";
    tmp(78047) := x"0021";
    tmp(78048) := x"0020";
    tmp(78049) := x"0800";
    tmp(78050) := x"0800";
    tmp(78051) := x"0800";
    tmp(78052) := x"1000";
    tmp(78053) := x"1000";
    tmp(78054) := x"1000";
    tmp(78055) := x"1000";
    tmp(78056) := x"1000";
    tmp(78057) := x"1020";
    tmp(78058) := x"1020";
    tmp(78059) := x"0800";
    tmp(78060) := x"0800";
    tmp(78061) := x"0800";
    tmp(78062) := x"1000";
    tmp(78063) := x"1000";
    tmp(78064) := x"1000";
    tmp(78065) := x"1000";
    tmp(78066) := x"1000";
    tmp(78067) := x"1000";
    tmp(78068) := x"1000";
    tmp(78069) := x"1000";
    tmp(78070) := x"1000";
    tmp(78071) := x"1000";
    tmp(78072) := x"1000";
    tmp(78073) := x"1000";
    tmp(78074) := x"1800";
    tmp(78075) := x"1800";
    tmp(78076) := x"1800";
    tmp(78077) := x"1800";
    tmp(78078) := x"1800";
    tmp(78079) := x"1000";
    tmp(78080) := x"1800";
    tmp(78081) := x"1800";
    tmp(78082) := x"1000";
    tmp(78083) := x"1000";
    tmp(78084) := x"1000";
    tmp(78085) := x"0800";
    tmp(78086) := x"0800";
    tmp(78087) := x"0800";
    tmp(78088) := x"0800";
    tmp(78089) := x"1000";
    tmp(78090) := x"1000";
    tmp(78091) := x"0800";
    tmp(78092) := x"0800";
    tmp(78093) := x"1000";
    tmp(78094) := x"1000";
    tmp(78095) := x"0800";
    tmp(78096) := x"0800";
    tmp(78097) := x"0800";
    tmp(78098) := x"0800";
    tmp(78099) := x"0800";
    tmp(78100) := x"0800";
    tmp(78101) := x"1000";
    tmp(78102) := x"0800";
    tmp(78103) := x"0800";
    tmp(78104) := x"0820";
    tmp(78105) := x"0020";
    tmp(78106) := x"0020";
    tmp(78107) := x"0020";
    tmp(78108) := x"0020";
    tmp(78109) := x"0020";
    tmp(78110) := x"0020";
    tmp(78111) := x"0000";
    tmp(78112) := x"0000";
    tmp(78113) := x"0000";
    tmp(78114) := x"0000";
    tmp(78115) := x"0000";
    tmp(78116) := x"0000";
    tmp(78117) := x"0000";
    tmp(78118) := x"0000";
    tmp(78119) := x"0000";
    tmp(78120) := x"0000";
    tmp(78121) := x"0000";
    tmp(78122) := x"0000";
    tmp(78123) := x"0000";
    tmp(78124) := x"0000";
    tmp(78125) := x"0000";
    tmp(78126) := x"0000";
    tmp(78127) := x"0000";
    tmp(78128) := x"0000";
    tmp(78129) := x"0000";
    tmp(78130) := x"0000";
    tmp(78131) := x"0000";
    tmp(78132) := x"0000";
    tmp(78133) := x"0000";
    tmp(78134) := x"0000";
    tmp(78135) := x"0000";
    tmp(78136) := x"0000";
    tmp(78137) := x"0000";
    tmp(78138) := x"0000";
    tmp(78139) := x"0000";
    tmp(78140) := x"0000";
    tmp(78141) := x"0000";
    tmp(78142) := x"0000";
    tmp(78143) := x"0000";
    tmp(78144) := x"0000";
    tmp(78145) := x"0000";
    tmp(78146) := x"0000";
    tmp(78147) := x"0000";
    tmp(78148) := x"0000";
    tmp(78149) := x"0000";
    tmp(78150) := x"0000";
    tmp(78151) := x"0000";
    tmp(78152) := x"0000";
    tmp(78153) := x"0000";
    tmp(78154) := x"0000";
    tmp(78155) := x"0000";
    tmp(78156) := x"0000";
    tmp(78157) := x"0000";
    tmp(78158) := x"0000";
    tmp(78159) := x"0000";
    tmp(78160) := x"0000";
    tmp(78161) := x"0000";
    tmp(78162) := x"0000";
    tmp(78163) := x"0000";
    tmp(78164) := x"0000";
    tmp(78165) := x"0000";
    tmp(78166) := x"0000";
    tmp(78167) := x"0000";
    tmp(78168) := x"0000";
    tmp(78169) := x"0000";
    tmp(78170) := x"0000";
    tmp(78171) := x"0000";
    tmp(78172) := x"0000";
    tmp(78173) := x"0000";
    tmp(78174) := x"0000";
    tmp(78175) := x"0000";
    tmp(78176) := x"0000";
    tmp(78177) := x"0000";
    tmp(78178) := x"0000";
    tmp(78179) := x"0000";
    tmp(78180) := x"0000";
    tmp(78181) := x"0000";
    tmp(78182) := x"0000";
    tmp(78183) := x"0000";
    tmp(78184) := x"0000";
    tmp(78185) := x"0000";
    tmp(78186) := x"0000";
    tmp(78187) := x"0000";
    tmp(78188) := x"0000";
    tmp(78189) := x"0000";
    tmp(78190) := x"0000";
    tmp(78191) := x"0000";
    tmp(78192) := x"0000";
    tmp(78193) := x"0000";
    tmp(78194) := x"0000";
    tmp(78195) := x"0000";
    tmp(78196) := x"0000";
    tmp(78197) := x"0000";
    tmp(78198) := x"0000";
    tmp(78199) := x"0000";
    tmp(78200) := x"0000";
    tmp(78201) := x"0000";
    tmp(78202) := x"0000";
    tmp(78203) := x"0000";
    tmp(78204) := x"0000";
    tmp(78205) := x"0000";
    tmp(78206) := x"0000";
    tmp(78207) := x"0000";
    tmp(78208) := x"0000";
    tmp(78209) := x"0000";
    tmp(78210) := x"0000";
    tmp(78211) := x"0000";
    tmp(78212) := x"0000";
    tmp(78213) := x"0000";
    tmp(78214) := x"0000";
    tmp(78215) := x"0000";
    tmp(78216) := x"0000";
    tmp(78217) := x"0000";
    tmp(78218) := x"0000";
    tmp(78219) := x"0000";
    tmp(78220) := x"0000";
    tmp(78221) := x"0000";
    tmp(78222) := x"0000";
    tmp(78223) := x"0000";
    tmp(78224) := x"0000";
    tmp(78225) := x"0000";
    tmp(78226) := x"0000";
    tmp(78227) := x"0000";
    tmp(78228) := x"0000";
    tmp(78229) := x"0000";
    tmp(78230) := x"0000";
    tmp(78231) := x"0000";
    tmp(78232) := x"0000";
    tmp(78233) := x"0000";
    tmp(78234) := x"0000";
    tmp(78235) := x"0000";
    tmp(78236) := x"0000";
    tmp(78237) := x"0000";
    tmp(78238) := x"0000";
    tmp(78239) := x"0000";
    tmp(78240) := x"0000";
    tmp(78241) := x"0020";
    tmp(78242) := x"0020";
    tmp(78243) := x"0020";
    tmp(78244) := x"0000";
    tmp(78245) := x"0000";
    tmp(78246) := x"0000";
    tmp(78247) := x"0020";
    tmp(78248) := x"0020";
    tmp(78249) := x"0020";
    tmp(78250) := x"0020";
    tmp(78251) := x"0020";
    tmp(78252) := x"0020";
    tmp(78253) := x"0020";
    tmp(78254) := x"0040";
    tmp(78255) := x"0040";
    tmp(78256) := x"0040";
    tmp(78257) := x"0040";
    tmp(78258) := x"0040";
    tmp(78259) := x"0040";
    tmp(78260) := x"0040";
    tmp(78261) := x"0040";
    tmp(78262) := x"0040";
    tmp(78263) := x"0040";
    tmp(78264) := x"0040";
    tmp(78265) := x"0040";
    tmp(78266) := x"0040";
    tmp(78267) := x"0040";
    tmp(78268) := x"0040";
    tmp(78269) := x"0040";
    tmp(78270) := x"0040";
    tmp(78271) := x"0040";
    tmp(78272) := x"0040";
    tmp(78273) := x"0040";
    tmp(78274) := x"0040";
    tmp(78275) := x"0040";
    tmp(78276) := x"0040";
    tmp(78277) := x"0040";
    tmp(78278) := x"0040";
    tmp(78279) := x"0040";
    tmp(78280) := x"0041";
    tmp(78281) := x"0041";
    tmp(78282) := x"0041";
    tmp(78283) := x"0041";
    tmp(78284) := x"0041";
    tmp(78285) := x"0021";
    tmp(78286) := x"0021";
    tmp(78287) := x"0021";
    tmp(78288) := x"0020";
    tmp(78289) := x"0820";
    tmp(78290) := x"0800";
    tmp(78291) := x"0800";
    tmp(78292) := x"1000";
    tmp(78293) := x"1000";
    tmp(78294) := x"1000";
    tmp(78295) := x"1000";
    tmp(78296) := x"1000";
    tmp(78297) := x"1000";
    tmp(78298) := x"1000";
    tmp(78299) := x"1000";
    tmp(78300) := x"0800";
    tmp(78301) := x"0800";
    tmp(78302) := x"1000";
    tmp(78303) := x"1000";
    tmp(78304) := x"1000";
    tmp(78305) := x"1000";
    tmp(78306) := x"1000";
    tmp(78307) := x"1000";
    tmp(78308) := x"1000";
    tmp(78309) := x"1000";
    tmp(78310) := x"1000";
    tmp(78311) := x"1800";
    tmp(78312) := x"1800";
    tmp(78313) := x"1800";
    tmp(78314) := x"1800";
    tmp(78315) := x"1000";
    tmp(78316) := x"1000";
    tmp(78317) := x"1800";
    tmp(78318) := x"1000";
    tmp(78319) := x"1000";
    tmp(78320) := x"1000";
    tmp(78321) := x"1000";
    tmp(78322) := x"0800";
    tmp(78323) := x"0800";
    tmp(78324) := x"0000";
    tmp(78325) := x"0800";
    tmp(78326) := x"0800";
    tmp(78327) := x"1000";
    tmp(78328) := x"1000";
    tmp(78329) := x"1000";
    tmp(78330) := x"1000";
    tmp(78331) := x"0800";
    tmp(78332) := x"0000";
    tmp(78333) := x"0800";
    tmp(78334) := x"1000";
    tmp(78335) := x"1820";
    tmp(78336) := x"0800";
    tmp(78337) := x"0000";
    tmp(78338) := x"0000";
    tmp(78339) := x"0800";
    tmp(78340) := x"1000";
    tmp(78341) := x"1800";
    tmp(78342) := x"1020";
    tmp(78343) := x"0820";
    tmp(78344) := x"0000";
    tmp(78345) := x"0020";
    tmp(78346) := x"0020";
    tmp(78347) := x"0020";
    tmp(78348) := x"0020";
    tmp(78349) := x"0020";
    tmp(78350) := x"0020";
    tmp(78351) := x"0000";
    tmp(78352) := x"0000";
    tmp(78353) := x"0000";
    tmp(78354) := x"0000";
    tmp(78355) := x"0000";
    tmp(78356) := x"0000";
    tmp(78357) := x"0000";
    tmp(78358) := x"0000";
    tmp(78359) := x"0000";
    tmp(78360) := x"0000";
    tmp(78361) := x"0000";
    tmp(78362) := x"0000";
    tmp(78363) := x"0000";
    tmp(78364) := x"0000";
    tmp(78365) := x"0000";
    tmp(78366) := x"0000";
    tmp(78367) := x"0000";
    tmp(78368) := x"0000";
    tmp(78369) := x"0000";
    tmp(78370) := x"0000";
    tmp(78371) := x"0000";
    tmp(78372) := x"0000";
    tmp(78373) := x"0000";
    tmp(78374) := x"0000";
    tmp(78375) := x"0000";
    tmp(78376) := x"0000";
    tmp(78377) := x"0000";
    tmp(78378) := x"0000";
    tmp(78379) := x"0000";
    tmp(78380) := x"0000";
    tmp(78381) := x"0000";
    tmp(78382) := x"0000";
    tmp(78383) := x"0000";
    tmp(78384) := x"0000";
    tmp(78385) := x"0000";
    tmp(78386) := x"0000";
    tmp(78387) := x"0000";
    tmp(78388) := x"0000";
    tmp(78389) := x"0000";
    tmp(78390) := x"0000";
    tmp(78391) := x"0000";
    tmp(78392) := x"0000";
    tmp(78393) := x"0000";
    tmp(78394) := x"0000";
    tmp(78395) := x"0000";
    tmp(78396) := x"0000";
    tmp(78397) := x"0000";
    tmp(78398) := x"0000";
    tmp(78399) := x"0000";
    tmp(78400) := x"0000";
    tmp(78401) := x"0000";
    tmp(78402) := x"0000";
    tmp(78403) := x"0000";
    tmp(78404) := x"0000";
    tmp(78405) := x"0000";
    tmp(78406) := x"0000";
    tmp(78407) := x"0000";
    tmp(78408) := x"0000";
    tmp(78409) := x"0000";
    tmp(78410) := x"0000";
    tmp(78411) := x"0000";
    tmp(78412) := x"0000";
    tmp(78413) := x"0000";
    tmp(78414) := x"0000";
    tmp(78415) := x"0000";
    tmp(78416) := x"0000";
    tmp(78417) := x"0000";
    tmp(78418) := x"0000";
    tmp(78419) := x"0000";
    tmp(78420) := x"0000";
    tmp(78421) := x"0000";
    tmp(78422) := x"0000";
    tmp(78423) := x"0000";
    tmp(78424) := x"0000";
    tmp(78425) := x"0000";
    tmp(78426) := x"0000";
    tmp(78427) := x"0000";
    tmp(78428) := x"0000";
    tmp(78429) := x"0000";
    tmp(78430) := x"0000";
    tmp(78431) := x"0000";
    tmp(78432) := x"0000";
    tmp(78433) := x"0000";
    tmp(78434) := x"0000";
    tmp(78435) := x"0000";
    tmp(78436) := x"0000";
    tmp(78437) := x"0000";
    tmp(78438) := x"0000";
    tmp(78439) := x"0000";
    tmp(78440) := x"0000";
    tmp(78441) := x"0000";
    tmp(78442) := x"0000";
    tmp(78443) := x"0000";
    tmp(78444) := x"0000";
    tmp(78445) := x"0000";
    tmp(78446) := x"0000";
    tmp(78447) := x"0000";
    tmp(78448) := x"0000";
    tmp(78449) := x"0000";
    tmp(78450) := x"0000";
    tmp(78451) := x"0000";
    tmp(78452) := x"0000";
    tmp(78453) := x"0000";
    tmp(78454) := x"0000";
    tmp(78455) := x"0000";
    tmp(78456) := x"0000";
    tmp(78457) := x"0000";
    tmp(78458) := x"0000";
    tmp(78459) := x"0000";
    tmp(78460) := x"0000";
    tmp(78461) := x"0000";
    tmp(78462) := x"0000";
    tmp(78463) := x"0000";
    tmp(78464) := x"0000";
    tmp(78465) := x"0000";
    tmp(78466) := x"0000";
    tmp(78467) := x"0000";
    tmp(78468) := x"0000";
    tmp(78469) := x"0000";
    tmp(78470) := x"0000";
    tmp(78471) := x"0000";
    tmp(78472) := x"0000";
    tmp(78473) := x"0000";
    tmp(78474) := x"0000";
    tmp(78475) := x"0000";
    tmp(78476) := x"0000";
    tmp(78477) := x"0000";
    tmp(78478) := x"0000";
    tmp(78479) := x"0000";
    tmp(78480) := x"0000";
    tmp(78481) := x"0020";
    tmp(78482) := x"0020";
    tmp(78483) := x"0020";
    tmp(78484) := x"0020";
    tmp(78485) := x"0000";
    tmp(78486) := x"0000";
    tmp(78487) := x"0000";
    tmp(78488) := x"0020";
    tmp(78489) := x"0020";
    tmp(78490) := x"0020";
    tmp(78491) := x"0020";
    tmp(78492) := x"0020";
    tmp(78493) := x"0020";
    tmp(78494) := x"0020";
    tmp(78495) := x"0020";
    tmp(78496) := x"0020";
    tmp(78497) := x"0020";
    tmp(78498) := x"0040";
    tmp(78499) := x"0040";
    tmp(78500) := x"0040";
    tmp(78501) := x"0040";
    tmp(78502) := x"0040";
    tmp(78503) := x"0040";
    tmp(78504) := x"0040";
    tmp(78505) := x"0040";
    tmp(78506) := x"0040";
    tmp(78507) := x"0040";
    tmp(78508) := x"0040";
    tmp(78509) := x"0040";
    tmp(78510) := x"0040";
    tmp(78511) := x"0040";
    tmp(78512) := x"0040";
    tmp(78513) := x"0040";
    tmp(78514) := x"0040";
    tmp(78515) := x"0040";
    tmp(78516) := x"0040";
    tmp(78517) := x"0040";
    tmp(78518) := x"0040";
    tmp(78519) := x"0041";
    tmp(78520) := x"0041";
    tmp(78521) := x"0041";
    tmp(78522) := x"0041";
    tmp(78523) := x"0041";
    tmp(78524) := x"0041";
    tmp(78525) := x"0041";
    tmp(78526) := x"0021";
    tmp(78527) := x"0021";
    tmp(78528) := x"0021";
    tmp(78529) := x"0020";
    tmp(78530) := x"0020";
    tmp(78531) := x"0800";
    tmp(78532) := x"0800";
    tmp(78533) := x"1000";
    tmp(78534) := x"1000";
    tmp(78535) := x"1800";
    tmp(78536) := x"1800";
    tmp(78537) := x"1800";
    tmp(78538) := x"1000";
    tmp(78539) := x"1000";
    tmp(78540) := x"0800";
    tmp(78541) := x"0800";
    tmp(78542) := x"1000";
    tmp(78543) := x"1000";
    tmp(78544) := x"1000";
    tmp(78545) := x"1000";
    tmp(78546) := x"1800";
    tmp(78547) := x"1800";
    tmp(78548) := x"2000";
    tmp(78549) := x"2020";
    tmp(78550) := x"2020";
    tmp(78551) := x"2000";
    tmp(78552) := x"2000";
    tmp(78553) := x"1800";
    tmp(78554) := x"1000";
    tmp(78555) := x"1000";
    tmp(78556) := x"1800";
    tmp(78557) := x"1000";
    tmp(78558) := x"1000";
    tmp(78559) := x"1000";
    tmp(78560) := x"1000";
    tmp(78561) := x"0800";
    tmp(78562) := x"0800";
    tmp(78563) := x"0800";
    tmp(78564) := x"0800";
    tmp(78565) := x"1000";
    tmp(78566) := x"1020";
    tmp(78567) := x"1020";
    tmp(78568) := x"0800";
    tmp(78569) := x"0000";
    tmp(78570) := x"0000";
    tmp(78571) := x"0000";
    tmp(78572) := x"0800";
    tmp(78573) := x"2020";
    tmp(78574) := x"1820";
    tmp(78575) := x"0800";
    tmp(78576) := x"0000";
    tmp(78577) := x"0000";
    tmp(78578) := x"0800";
    tmp(78579) := x"1000";
    tmp(78580) := x"1800";
    tmp(78581) := x"1820";
    tmp(78582) := x"0820";
    tmp(78583) := x"0000";
    tmp(78584) := x"0000";
    tmp(78585) := x"0000";
    tmp(78586) := x"0020";
    tmp(78587) := x"0020";
    tmp(78588) := x"0020";
    tmp(78589) := x"0020";
    tmp(78590) := x"0020";
    tmp(78591) := x"0000";
    tmp(78592) := x"0000";
    tmp(78593) := x"0000";
    tmp(78594) := x"0000";
    tmp(78595) := x"0000";
    tmp(78596) := x"0000";
    tmp(78597) := x"0000";
    tmp(78598) := x"0000";
    tmp(78599) := x"0000";
    tmp(78600) := x"0000";
    tmp(78601) := x"0000";
    tmp(78602) := x"0000";
    tmp(78603) := x"0000";
    tmp(78604) := x"0000";
    tmp(78605) := x"0000";
    tmp(78606) := x"0000";
    tmp(78607) := x"0000";
    tmp(78608) := x"0000";
    tmp(78609) := x"0000";
    tmp(78610) := x"0000";
    tmp(78611) := x"0000";
    tmp(78612) := x"0000";
    tmp(78613) := x"0000";
    tmp(78614) := x"0000";
    tmp(78615) := x"0000";
    tmp(78616) := x"0000";
    tmp(78617) := x"0000";
    tmp(78618) := x"0000";
    tmp(78619) := x"0000";
    tmp(78620) := x"0000";
    tmp(78621) := x"0000";
    tmp(78622) := x"0000";
    tmp(78623) := x"0000";
    tmp(78624) := x"0000";
    tmp(78625) := x"0000";
    tmp(78626) := x"0000";
    tmp(78627) := x"0000";
    tmp(78628) := x"0000";
    tmp(78629) := x"0000";
    tmp(78630) := x"0000";
    tmp(78631) := x"0000";
    tmp(78632) := x"0000";
    tmp(78633) := x"0000";
    tmp(78634) := x"0000";
    tmp(78635) := x"0000";
    tmp(78636) := x"0000";
    tmp(78637) := x"0000";
    tmp(78638) := x"0000";
    tmp(78639) := x"0000";
    tmp(78640) := x"0000";
    tmp(78641) := x"0000";
    tmp(78642) := x"0000";
    tmp(78643) := x"0000";
    tmp(78644) := x"0000";
    tmp(78645) := x"0000";
    tmp(78646) := x"0000";
    tmp(78647) := x"0000";
    tmp(78648) := x"0000";
    tmp(78649) := x"0000";
    tmp(78650) := x"0000";
    tmp(78651) := x"0000";
    tmp(78652) := x"0000";
    tmp(78653) := x"0000";
    tmp(78654) := x"0000";
    tmp(78655) := x"0000";
    tmp(78656) := x"0000";
    tmp(78657) := x"0000";
    tmp(78658) := x"0000";
    tmp(78659) := x"0000";
    tmp(78660) := x"0000";
    tmp(78661) := x"0000";
    tmp(78662) := x"0000";
    tmp(78663) := x"0000";
    tmp(78664) := x"0000";
    tmp(78665) := x"0000";
    tmp(78666) := x"0000";
    tmp(78667) := x"0000";
    tmp(78668) := x"0000";
    tmp(78669) := x"0000";
    tmp(78670) := x"0000";
    tmp(78671) := x"0000";
    tmp(78672) := x"0000";
    tmp(78673) := x"0000";
    tmp(78674) := x"0000";
    tmp(78675) := x"0000";
    tmp(78676) := x"0000";
    tmp(78677) := x"0000";
    tmp(78678) := x"0000";
    tmp(78679) := x"0000";
    tmp(78680) := x"0000";
    tmp(78681) := x"0000";
    tmp(78682) := x"0000";
    tmp(78683) := x"0000";
    tmp(78684) := x"0000";
    tmp(78685) := x"0000";
    tmp(78686) := x"0000";
    tmp(78687) := x"0000";
    tmp(78688) := x"0000";
    tmp(78689) := x"0000";
    tmp(78690) := x"0000";
    tmp(78691) := x"0000";
    tmp(78692) := x"0000";
    tmp(78693) := x"0000";
    tmp(78694) := x"0000";
    tmp(78695) := x"0000";
    tmp(78696) := x"0000";
    tmp(78697) := x"0000";
    tmp(78698) := x"0000";
    tmp(78699) := x"0000";
    tmp(78700) := x"0000";
    tmp(78701) := x"0000";
    tmp(78702) := x"0000";
    tmp(78703) := x"0000";
    tmp(78704) := x"0000";
    tmp(78705) := x"0000";
    tmp(78706) := x"0000";
    tmp(78707) := x"0000";
    tmp(78708) := x"0000";
    tmp(78709) := x"0000";
    tmp(78710) := x"0000";
    tmp(78711) := x"0000";
    tmp(78712) := x"0000";
    tmp(78713) := x"0000";
    tmp(78714) := x"0000";
    tmp(78715) := x"0000";
    tmp(78716) := x"0000";
    tmp(78717) := x"0000";
    tmp(78718) := x"0000";
    tmp(78719) := x"0000";
    tmp(78720) := x"0000";
    tmp(78721) := x"0020";
    tmp(78722) := x"0020";
    tmp(78723) := x"0020";
    tmp(78724) := x"0020";
    tmp(78725) := x"0020";
    tmp(78726) := x"0020";
    tmp(78727) := x"0020";
    tmp(78728) := x"0000";
    tmp(78729) := x"0020";
    tmp(78730) := x"0020";
    tmp(78731) := x"0020";
    tmp(78732) := x"0020";
    tmp(78733) := x"0020";
    tmp(78734) := x"0020";
    tmp(78735) := x"0020";
    tmp(78736) := x"0020";
    tmp(78737) := x"0020";
    tmp(78738) := x"0020";
    tmp(78739) := x"0020";
    tmp(78740) := x"0020";
    tmp(78741) := x"0040";
    tmp(78742) := x"0040";
    tmp(78743) := x"0040";
    tmp(78744) := x"0040";
    tmp(78745) := x"0040";
    tmp(78746) := x"0040";
    tmp(78747) := x"0040";
    tmp(78748) := x"0040";
    tmp(78749) := x"0040";
    tmp(78750) := x"0040";
    tmp(78751) := x"0040";
    tmp(78752) := x"0040";
    tmp(78753) := x"0040";
    tmp(78754) := x"0040";
    tmp(78755) := x"0040";
    tmp(78756) := x"0040";
    tmp(78757) := x"0040";
    tmp(78758) := x"0040";
    tmp(78759) := x"0040";
    tmp(78760) := x"0041";
    tmp(78761) := x"0041";
    tmp(78762) := x"0041";
    tmp(78763) := x"0041";
    tmp(78764) := x"0041";
    tmp(78765) := x"0041";
    tmp(78766) := x"0041";
    tmp(78767) := x"0041";
    tmp(78768) := x"0021";
    tmp(78769) := x"0021";
    tmp(78770) := x"0020";
    tmp(78771) := x"0020";
    tmp(78772) := x"0000";
    tmp(78773) := x"0800";
    tmp(78774) := x"1000";
    tmp(78775) := x"1000";
    tmp(78776) := x"1800";
    tmp(78777) := x"1800";
    tmp(78778) := x"1000";
    tmp(78779) := x"0800";
    tmp(78780) := x"0800";
    tmp(78781) := x"1000";
    tmp(78782) := x"1000";
    tmp(78783) := x"1000";
    tmp(78784) := x"1800";
    tmp(78785) := x"1800";
    tmp(78786) := x"1800";
    tmp(78787) := x"1800";
    tmp(78788) := x"1800";
    tmp(78789) := x"1800";
    tmp(78790) := x"1800";
    tmp(78791) := x"2020";
    tmp(78792) := x"1820";
    tmp(78793) := x"1000";
    tmp(78794) := x"1000";
    tmp(78795) := x"1000";
    tmp(78796) := x"1000";
    tmp(78797) := x"1000";
    tmp(78798) := x"1000";
    tmp(78799) := x"1000";
    tmp(78800) := x"1000";
    tmp(78801) := x"0800";
    tmp(78802) := x"0800";
    tmp(78803) := x"1000";
    tmp(78804) := x"1000";
    tmp(78805) := x"1000";
    tmp(78806) := x"0800";
    tmp(78807) := x"0000";
    tmp(78808) := x"0000";
    tmp(78809) := x"0000";
    tmp(78810) := x"0000";
    tmp(78811) := x"0000";
    tmp(78812) := x"2020";
    tmp(78813) := x"1000";
    tmp(78814) := x"0800";
    tmp(78815) := x"0000";
    tmp(78816) := x"0800";
    tmp(78817) := x"0800";
    tmp(78818) := x"1800";
    tmp(78819) := x"1800";
    tmp(78820) := x"1820";
    tmp(78821) := x"0820";
    tmp(78822) := x"0000";
    tmp(78823) := x"0000";
    tmp(78824) := x"0000";
    tmp(78825) := x"0000";
    tmp(78826) := x"0000";
    tmp(78827) := x"0000";
    tmp(78828) := x"0000";
    tmp(78829) := x"0000";
    tmp(78830) := x"0000";
    tmp(78831) := x"0000";
    tmp(78832) := x"0000";
    tmp(78833) := x"0000";
    tmp(78834) := x"0000";
    tmp(78835) := x"0000";
    tmp(78836) := x"0000";
    tmp(78837) := x"0000";
    tmp(78838) := x"0000";
    tmp(78839) := x"0000";
    tmp(78840) := x"0000";
    tmp(78841) := x"0000";
    tmp(78842) := x"0000";
    tmp(78843) := x"0000";
    tmp(78844) := x"0000";
    tmp(78845) := x"0000";
    tmp(78846) := x"0000";
    tmp(78847) := x"0000";
    tmp(78848) := x"0000";
    tmp(78849) := x"0000";
    tmp(78850) := x"0000";
    tmp(78851) := x"0000";
    tmp(78852) := x"0000";
    tmp(78853) := x"0000";
    tmp(78854) := x"0000";
    tmp(78855) := x"0000";
    tmp(78856) := x"0000";
    tmp(78857) := x"0000";
    tmp(78858) := x"0000";
    tmp(78859) := x"0000";
    tmp(78860) := x"0000";
    tmp(78861) := x"0000";
    tmp(78862) := x"0000";
    tmp(78863) := x"0000";
    tmp(78864) := x"0000";
    tmp(78865) := x"0000";
    tmp(78866) := x"0000";
    tmp(78867) := x"0000";
    tmp(78868) := x"0000";
    tmp(78869) := x"0000";
    tmp(78870) := x"0000";
    tmp(78871) := x"0000";
    tmp(78872) := x"0000";
    tmp(78873) := x"0000";
    tmp(78874) := x"0000";
    tmp(78875) := x"0000";
    tmp(78876) := x"0000";
    tmp(78877) := x"0000";
    tmp(78878) := x"0000";
    tmp(78879) := x"0000";
    tmp(78880) := x"0000";
    tmp(78881) := x"0000";
    tmp(78882) := x"0000";
    tmp(78883) := x"0000";
    tmp(78884) := x"0000";
    tmp(78885) := x"0000";
    tmp(78886) := x"0000";
    tmp(78887) := x"0000";
    tmp(78888) := x"0000";
    tmp(78889) := x"0000";
    tmp(78890) := x"0000";
    tmp(78891) := x"0000";
    tmp(78892) := x"0000";
    tmp(78893) := x"0000";
    tmp(78894) := x"0000";
    tmp(78895) := x"0000";
    tmp(78896) := x"0000";
    tmp(78897) := x"0000";
    tmp(78898) := x"0000";
    tmp(78899) := x"0000";
    tmp(78900) := x"0000";
    tmp(78901) := x"0000";
    tmp(78902) := x"0000";
    tmp(78903) := x"0000";
    tmp(78904) := x"0000";
    tmp(78905) := x"0000";
    tmp(78906) := x"0000";
    tmp(78907) := x"0000";
    tmp(78908) := x"0000";
    tmp(78909) := x"0000";
    tmp(78910) := x"0000";
    tmp(78911) := x"0000";
    tmp(78912) := x"0000";
    tmp(78913) := x"0000";
    tmp(78914) := x"0000";
    tmp(78915) := x"0000";
    tmp(78916) := x"0000";
    tmp(78917) := x"0000";
    tmp(78918) := x"0000";
    tmp(78919) := x"0000";
    tmp(78920) := x"0000";
    tmp(78921) := x"0000";
    tmp(78922) := x"0000";
    tmp(78923) := x"0000";
    tmp(78924) := x"0000";
    tmp(78925) := x"0000";
    tmp(78926) := x"0000";
    tmp(78927) := x"0000";
    tmp(78928) := x"0000";
    tmp(78929) := x"0000";
    tmp(78930) := x"0000";
    tmp(78931) := x"0000";
    tmp(78932) := x"0000";
    tmp(78933) := x"0000";
    tmp(78934) := x"0000";
    tmp(78935) := x"0000";
    tmp(78936) := x"0000";
    tmp(78937) := x"0000";
    tmp(78938) := x"0000";
    tmp(78939) := x"0000";
    tmp(78940) := x"0000";
    tmp(78941) := x"0000";
    tmp(78942) := x"0000";
    tmp(78943) := x"0000";
    tmp(78944) := x"0000";
    tmp(78945) := x"0000";
    tmp(78946) := x"0000";
    tmp(78947) := x"0000";
    tmp(78948) := x"0000";
    tmp(78949) := x"0000";
    tmp(78950) := x"0000";
    tmp(78951) := x"0000";
    tmp(78952) := x"0000";
    tmp(78953) := x"0000";
    tmp(78954) := x"0000";
    tmp(78955) := x"0000";
    tmp(78956) := x"0000";
    tmp(78957) := x"0000";
    tmp(78958) := x"0000";
    tmp(78959) := x"0000";
    tmp(78960) := x"0000";
    tmp(78961) := x"0020";
    tmp(78962) := x"0020";
    tmp(78963) := x"0020";
    tmp(78964) := x"0020";
    tmp(78965) := x"0020";
    tmp(78966) := x"0020";
    tmp(78967) := x"0020";
    tmp(78968) := x"0020";
    tmp(78969) := x"0020";
    tmp(78970) := x"0020";
    tmp(78971) := x"0020";
    tmp(78972) := x"0020";
    tmp(78973) := x"0040";
    tmp(78974) := x"0040";
    tmp(78975) := x"0020";
    tmp(78976) := x"0020";
    tmp(78977) := x"0020";
    tmp(78978) := x"0020";
    tmp(78979) := x"0020";
    tmp(78980) := x"0020";
    tmp(78981) := x"0020";
    tmp(78982) := x"0020";
    tmp(78983) := x"0020";
    tmp(78984) := x"0020";
    tmp(78985) := x"0020";
    tmp(78986) := x"0040";
    tmp(78987) := x"0040";
    tmp(78988) := x"0040";
    tmp(78989) := x"0040";
    tmp(78990) := x"0040";
    tmp(78991) := x"0040";
    tmp(78992) := x"0040";
    tmp(78993) := x"0040";
    tmp(78994) := x"0040";
    tmp(78995) := x"0040";
    tmp(78996) := x"0040";
    tmp(78997) := x"0040";
    tmp(78998) := x"0040";
    tmp(78999) := x"0040";
    tmp(79000) := x"0040";
    tmp(79001) := x"0041";
    tmp(79002) := x"0041";
    tmp(79003) := x"0041";
    tmp(79004) := x"0041";
    tmp(79005) := x"0041";
    tmp(79006) := x"0041";
    tmp(79007) := x"0041";
    tmp(79008) := x"0041";
    tmp(79009) := x"0020";
    tmp(79010) := x"0020";
    tmp(79011) := x"0020";
    tmp(79012) := x"0020";
    tmp(79013) := x"0000";
    tmp(79014) := x"0800";
    tmp(79015) := x"0800";
    tmp(79016) := x"1000";
    tmp(79017) := x"1000";
    tmp(79018) := x"0800";
    tmp(79019) := x"0800";
    tmp(79020) := x"0800";
    tmp(79021) := x"0800";
    tmp(79022) := x"1000";
    tmp(79023) := x"1000";
    tmp(79024) := x"1000";
    tmp(79025) := x"1000";
    tmp(79026) := x"1000";
    tmp(79027) := x"1800";
    tmp(79028) := x"1800";
    tmp(79029) := x"1800";
    tmp(79030) := x"1820";
    tmp(79031) := x"1820";
    tmp(79032) := x"1020";
    tmp(79033) := x"0800";
    tmp(79034) := x"1000";
    tmp(79035) := x"1000";
    tmp(79036) := x"1000";
    tmp(79037) := x"1000";
    tmp(79038) := x"0800";
    tmp(79039) := x"0800";
    tmp(79040) := x"0800";
    tmp(79041) := x"0800";
    tmp(79042) := x"0800";
    tmp(79043) := x"0800";
    tmp(79044) := x"0800";
    tmp(79045) := x"0000";
    tmp(79046) := x"0000";
    tmp(79047) := x"0000";
    tmp(79048) := x"0000";
    tmp(79049) := x"0000";
    tmp(79050) := x"0800";
    tmp(79051) := x"1000";
    tmp(79052) := x"0800";
    tmp(79053) := x"0800";
    tmp(79054) := x"0800";
    tmp(79055) := x"0800";
    tmp(79056) := x"0800";
    tmp(79057) := x"1800";
    tmp(79058) := x"1800";
    tmp(79059) := x"1800";
    tmp(79060) := x"0820";
    tmp(79061) := x"0000";
    tmp(79062) := x"0000";
    tmp(79063) := x"0000";
    tmp(79064) := x"0000";
    tmp(79065) := x"0000";
    tmp(79066) := x"0000";
    tmp(79067) := x"0000";
    tmp(79068) := x"0000";
    tmp(79069) := x"0000";
    tmp(79070) := x"0000";
    tmp(79071) := x"0000";
    tmp(79072) := x"0000";
    tmp(79073) := x"0000";
    tmp(79074) := x"0000";
    tmp(79075) := x"0000";
    tmp(79076) := x"0000";
    tmp(79077) := x"0000";
    tmp(79078) := x"0000";
    tmp(79079) := x"0000";
    tmp(79080) := x"0000";
    tmp(79081) := x"0000";
    tmp(79082) := x"0000";
    tmp(79083) := x"0000";
    tmp(79084) := x"0000";
    tmp(79085) := x"0000";
    tmp(79086) := x"0000";
    tmp(79087) := x"0000";
    tmp(79088) := x"0000";
    tmp(79089) := x"0000";
    tmp(79090) := x"0000";
    tmp(79091) := x"0000";
    tmp(79092) := x"0000";
    tmp(79093) := x"0000";
    tmp(79094) := x"0000";
    tmp(79095) := x"0000";
    tmp(79096) := x"0000";
    tmp(79097) := x"0000";
    tmp(79098) := x"0000";
    tmp(79099) := x"0000";
    tmp(79100) := x"0000";
    tmp(79101) := x"0000";
    tmp(79102) := x"0000";
    tmp(79103) := x"0000";
    tmp(79104) := x"0000";
    tmp(79105) := x"0000";
    tmp(79106) := x"0000";
    tmp(79107) := x"0000";
    tmp(79108) := x"0000";
    tmp(79109) := x"0000";
    tmp(79110) := x"0000";
    tmp(79111) := x"0000";
    tmp(79112) := x"0000";
    tmp(79113) := x"0000";
    tmp(79114) := x"0000";
    tmp(79115) := x"0000";
    tmp(79116) := x"0000";
    tmp(79117) := x"0000";
    tmp(79118) := x"0000";
    tmp(79119) := x"0000";
    tmp(79120) := x"0000";
    tmp(79121) := x"0000";
    tmp(79122) := x"0000";
    tmp(79123) := x"0000";
    tmp(79124) := x"0000";
    tmp(79125) := x"0000";
    tmp(79126) := x"0000";
    tmp(79127) := x"0000";
    tmp(79128) := x"0000";
    tmp(79129) := x"0000";
    tmp(79130) := x"0000";
    tmp(79131) := x"0000";
    tmp(79132) := x"0000";
    tmp(79133) := x"0000";
    tmp(79134) := x"0000";
    tmp(79135) := x"0000";
    tmp(79136) := x"0000";
    tmp(79137) := x"0000";
    tmp(79138) := x"0000";
    tmp(79139) := x"0000";
    tmp(79140) := x"0000";
    tmp(79141) := x"0000";
    tmp(79142) := x"0000";
    tmp(79143) := x"0000";
    tmp(79144) := x"0000";
    tmp(79145) := x"0000";
    tmp(79146) := x"0000";
    tmp(79147) := x"0000";
    tmp(79148) := x"0000";
    tmp(79149) := x"0000";
    tmp(79150) := x"0000";
    tmp(79151) := x"0000";
    tmp(79152) := x"0000";
    tmp(79153) := x"0000";
    tmp(79154) := x"0000";
    tmp(79155) := x"0000";
    tmp(79156) := x"0000";
    tmp(79157) := x"0000";
    tmp(79158) := x"0000";
    tmp(79159) := x"0000";
    tmp(79160) := x"0000";
    tmp(79161) := x"0000";
    tmp(79162) := x"0000";
    tmp(79163) := x"0000";
    tmp(79164) := x"0000";
    tmp(79165) := x"0000";
    tmp(79166) := x"0000";
    tmp(79167) := x"0000";
    tmp(79168) := x"0000";
    tmp(79169) := x"0000";
    tmp(79170) := x"0000";
    tmp(79171) := x"0000";
    tmp(79172) := x"0000";
    tmp(79173) := x"0000";
    tmp(79174) := x"0000";
    tmp(79175) := x"0000";
    tmp(79176) := x"0000";
    tmp(79177) := x"0000";
    tmp(79178) := x"0000";
    tmp(79179) := x"0000";
    tmp(79180) := x"0000";
    tmp(79181) := x"0000";
    tmp(79182) := x"0000";
    tmp(79183) := x"0000";
    tmp(79184) := x"0000";
    tmp(79185) := x"0000";
    tmp(79186) := x"0000";
    tmp(79187) := x"0000";
    tmp(79188) := x"0000";
    tmp(79189) := x"0000";
    tmp(79190) := x"0000";
    tmp(79191) := x"0000";
    tmp(79192) := x"0000";
    tmp(79193) := x"0000";
    tmp(79194) := x"0000";
    tmp(79195) := x"0000";
    tmp(79196) := x"0000";
    tmp(79197) := x"0000";
    tmp(79198) := x"0000";
    tmp(79199) := x"0000";
    tmp(79200) := x"0000";
    tmp(79201) := x"0020";
    tmp(79202) := x"0020";
    tmp(79203) := x"0020";
    tmp(79204) := x"0020";
    tmp(79205) := x"0020";
    tmp(79206) := x"0020";
    tmp(79207) := x"0020";
    tmp(79208) := x"0020";
    tmp(79209) := x"0020";
    tmp(79210) := x"0020";
    tmp(79211) := x"0020";
    tmp(79212) := x"0020";
    tmp(79213) := x"0020";
    tmp(79214) := x"0020";
    tmp(79215) := x"0040";
    tmp(79216) := x"0040";
    tmp(79217) := x"0020";
    tmp(79218) := x"0020";
    tmp(79219) := x"0020";
    tmp(79220) := x"0020";
    tmp(79221) := x"0020";
    tmp(79222) := x"0020";
    tmp(79223) := x"0020";
    tmp(79224) := x"0020";
    tmp(79225) := x"0020";
    tmp(79226) := x"0020";
    tmp(79227) := x"0020";
    tmp(79228) := x"0020";
    tmp(79229) := x"0020";
    tmp(79230) := x"0020";
    tmp(79231) := x"0020";
    tmp(79232) := x"0020";
    tmp(79233) := x"0040";
    tmp(79234) := x"0040";
    tmp(79235) := x"0040";
    tmp(79236) := x"0040";
    tmp(79237) := x"0040";
    tmp(79238) := x"0040";
    tmp(79239) := x"0840";
    tmp(79240) := x"0840";
    tmp(79241) := x"0040";
    tmp(79242) := x"0040";
    tmp(79243) := x"0840";
    tmp(79244) := x"0840";
    tmp(79245) := x"0840";
    tmp(79246) := x"0840";
    tmp(79247) := x"0840";
    tmp(79248) := x"0840";
    tmp(79249) := x"0840";
    tmp(79250) := x"0820";
    tmp(79251) := x"0820";
    tmp(79252) := x"0820";
    tmp(79253) := x"0800";
    tmp(79254) := x"0800";
    tmp(79255) := x"0800";
    tmp(79256) := x"1000";
    tmp(79257) := x"0800";
    tmp(79258) := x"0800";
    tmp(79259) := x"0800";
    tmp(79260) := x"0800";
    tmp(79261) := x"1000";
    tmp(79262) := x"1000";
    tmp(79263) := x"1000";
    tmp(79264) := x"1000";
    tmp(79265) := x"1000";
    tmp(79266) := x"1800";
    tmp(79267) := x"1800";
    tmp(79268) := x"1800";
    tmp(79269) := x"1820";
    tmp(79270) := x"1820";
    tmp(79271) := x"1000";
    tmp(79272) := x"1000";
    tmp(79273) := x"1000";
    tmp(79274) := x"1800";
    tmp(79275) := x"1800";
    tmp(79276) := x"1800";
    tmp(79277) := x"1020";
    tmp(79278) := x"1020";
    tmp(79279) := x"0800";
    tmp(79280) := x"0000";
    tmp(79281) := x"0000";
    tmp(79282) := x"0000";
    tmp(79283) := x"0000";
    tmp(79284) := x"0000";
    tmp(79285) := x"0000";
    tmp(79286) := x"0000";
    tmp(79287) := x"0000";
    tmp(79288) := x"0000";
    tmp(79289) := x"0800";
    tmp(79290) := x"0800";
    tmp(79291) := x"0800";
    tmp(79292) := x"0800";
    tmp(79293) := x"0800";
    tmp(79294) := x"1000";
    tmp(79295) := x"1000";
    tmp(79296) := x"1800";
    tmp(79297) := x"1800";
    tmp(79298) := x"1000";
    tmp(79299) := x"0820";
    tmp(79300) := x"0000";
    tmp(79301) := x"0000";
    tmp(79302) := x"0000";
    tmp(79303) := x"0000";
    tmp(79304) := x"0000";
    tmp(79305) := x"0000";
    tmp(79306) := x"0000";
    tmp(79307) := x"0000";
    tmp(79308) := x"0000";
    tmp(79309) := x"0000";
    tmp(79310) := x"0000";
    tmp(79311) := x"0000";
    tmp(79312) := x"0000";
    tmp(79313) := x"0000";
    tmp(79314) := x"0000";
    tmp(79315) := x"0000";
    tmp(79316) := x"0000";
    tmp(79317) := x"0000";
    tmp(79318) := x"0000";
    tmp(79319) := x"0000";
    tmp(79320) := x"0000";
    tmp(79321) := x"0000";
    tmp(79322) := x"0000";
    tmp(79323) := x"0000";
    tmp(79324) := x"0000";
    tmp(79325) := x"0000";
    tmp(79326) := x"0000";
    tmp(79327) := x"0000";
    tmp(79328) := x"0000";
    tmp(79329) := x"0000";
    tmp(79330) := x"0000";
    tmp(79331) := x"0000";
    tmp(79332) := x"0000";
    tmp(79333) := x"0000";
    tmp(79334) := x"0000";
    tmp(79335) := x"0000";
    tmp(79336) := x"0000";
    tmp(79337) := x"0000";
    tmp(79338) := x"0000";
    tmp(79339) := x"0000";
    tmp(79340) := x"0000";
    tmp(79341) := x"0000";
    tmp(79342) := x"0000";
    tmp(79343) := x"0000";
    tmp(79344) := x"0000";
    tmp(79345) := x"0000";
    tmp(79346) := x"0000";
    tmp(79347) := x"0000";
    tmp(79348) := x"0000";
    tmp(79349) := x"0000";
    tmp(79350) := x"0000";
    tmp(79351) := x"0000";
    tmp(79352) := x"0000";
    tmp(79353) := x"0000";
    tmp(79354) := x"0000";
    tmp(79355) := x"0000";
    tmp(79356) := x"0000";
    tmp(79357) := x"0000";
    tmp(79358) := x"0000";
    tmp(79359) := x"0000";
    tmp(79360) := x"0000";
    tmp(79361) := x"0000";
    tmp(79362) := x"0000";
    tmp(79363) := x"0000";
    tmp(79364) := x"0000";
    tmp(79365) := x"0000";
    tmp(79366) := x"0000";
    tmp(79367) := x"0000";
    tmp(79368) := x"0000";
    tmp(79369) := x"0000";
    tmp(79370) := x"0000";
    tmp(79371) := x"0000";
    tmp(79372) := x"0000";
    tmp(79373) := x"0000";
    tmp(79374) := x"0000";
    tmp(79375) := x"0000";
    tmp(79376) := x"0000";
    tmp(79377) := x"0000";
    tmp(79378) := x"0000";
    tmp(79379) := x"0000";
    tmp(79380) := x"0000";
    tmp(79381) := x"0000";
    tmp(79382) := x"0000";
    tmp(79383) := x"0000";
    tmp(79384) := x"0000";
    tmp(79385) := x"0000";
    tmp(79386) := x"0000";
    tmp(79387) := x"0000";
    tmp(79388) := x"0000";
    tmp(79389) := x"0000";
    tmp(79390) := x"0000";
    tmp(79391) := x"0000";
    tmp(79392) := x"0000";
    tmp(79393) := x"0000";
    tmp(79394) := x"0000";
    tmp(79395) := x"0000";
    tmp(79396) := x"0000";
    tmp(79397) := x"0000";
    tmp(79398) := x"0000";
    tmp(79399) := x"0000";
    tmp(79400) := x"0000";
    tmp(79401) := x"0000";
    tmp(79402) := x"0000";
    tmp(79403) := x"0000";
    tmp(79404) := x"0000";
    tmp(79405) := x"0000";
    tmp(79406) := x"0000";
    tmp(79407) := x"0000";
    tmp(79408) := x"0000";
    tmp(79409) := x"0000";
    tmp(79410) := x"0000";
    tmp(79411) := x"0000";
    tmp(79412) := x"0000";
    tmp(79413) := x"0000";
    tmp(79414) := x"0000";
    tmp(79415) := x"0000";
    tmp(79416) := x"0000";
    tmp(79417) := x"0000";
    tmp(79418) := x"0000";
    tmp(79419) := x"0000";
    tmp(79420) := x"0000";
    tmp(79421) := x"0000";
    tmp(79422) := x"0000";
    tmp(79423) := x"0000";
    tmp(79424) := x"0000";
    tmp(79425) := x"0000";
    tmp(79426) := x"0000";
    tmp(79427) := x"0000";
    tmp(79428) := x"0000";
    tmp(79429) := x"0000";
    tmp(79430) := x"0000";
    tmp(79431) := x"0000";
    tmp(79432) := x"0000";
    tmp(79433) := x"0000";
    tmp(79434) := x"0000";
    tmp(79435) := x"0000";
    tmp(79436) := x"0000";
    tmp(79437) := x"0000";
    tmp(79438) := x"0000";
    tmp(79439) := x"0000";
    tmp(79440) := x"0000";
    tmp(79441) := x"0020";
    tmp(79442) := x"0020";
    tmp(79443) := x"0020";
    tmp(79444) := x"0020";
    tmp(79445) := x"0020";
    tmp(79446) := x"0020";
    tmp(79447) := x"0020";
    tmp(79448) := x"0020";
    tmp(79449) := x"0020";
    tmp(79450) := x"0020";
    tmp(79451) := x"0020";
    tmp(79452) := x"0020";
    tmp(79453) := x"0020";
    tmp(79454) := x"0020";
    tmp(79455) := x"0020";
    tmp(79456) := x"0020";
    tmp(79457) := x"0040";
    tmp(79458) := x"0020";
    tmp(79459) := x"0020";
    tmp(79460) := x"0020";
    tmp(79461) := x"0020";
    tmp(79462) := x"0020";
    tmp(79463) := x"0020";
    tmp(79464) := x"0020";
    tmp(79465) := x"0020";
    tmp(79466) := x"0020";
    tmp(79467) := x"0020";
    tmp(79468) := x"0020";
    tmp(79469) := x"0020";
    tmp(79470) := x"0020";
    tmp(79471) := x"0020";
    tmp(79472) := x"0020";
    tmp(79473) := x"0020";
    tmp(79474) := x"0020";
    tmp(79475) := x"0020";
    tmp(79476) := x"0020";
    tmp(79477) := x"0020";
    tmp(79478) := x"0820";
    tmp(79479) := x"0820";
    tmp(79480) := x"0820";
    tmp(79481) := x"0820";
    tmp(79482) := x"0820";
    tmp(79483) := x"0820";
    tmp(79484) := x"0820";
    tmp(79485) := x"0820";
    tmp(79486) := x"0820";
    tmp(79487) := x"0820";
    tmp(79488) := x"0820";
    tmp(79489) := x"0820";
    tmp(79490) := x"0800";
    tmp(79491) := x"0800";
    tmp(79492) := x"0800";
    tmp(79493) := x"0800";
    tmp(79494) := x"1000";
    tmp(79495) := x"1000";
    tmp(79496) := x"1000";
    tmp(79497) := x"0800";
    tmp(79498) := x"0800";
    tmp(79499) := x"0800";
    tmp(79500) := x"0800";
    tmp(79501) := x"1000";
    tmp(79502) := x"1000";
    tmp(79503) := x"1000";
    tmp(79504) := x"1000";
    tmp(79505) := x"1000";
    tmp(79506) := x"1000";
    tmp(79507) := x"1800";
    tmp(79508) := x"1800";
    tmp(79509) := x"1800";
    tmp(79510) := x"1800";
    tmp(79511) := x"1000";
    tmp(79512) := x"1000";
    tmp(79513) := x"1820";
    tmp(79514) := x"1820";
    tmp(79515) := x"1820";
    tmp(79516) := x"1020";
    tmp(79517) := x"1000";
    tmp(79518) := x"0800";
    tmp(79519) := x"0000";
    tmp(79520) := x"0000";
    tmp(79521) := x"0000";
    tmp(79522) := x"0000";
    tmp(79523) := x"0000";
    tmp(79524) := x"0000";
    tmp(79525) := x"0000";
    tmp(79526) := x"0000";
    tmp(79527) := x"0800";
    tmp(79528) := x"0800";
    tmp(79529) := x"0800";
    tmp(79530) := x"0800";
    tmp(79531) := x"0800";
    tmp(79532) := x"0800";
    tmp(79533) := x"1000";
    tmp(79534) := x"1000";
    tmp(79535) := x"1000";
    tmp(79536) := x"1000";
    tmp(79537) := x"1000";
    tmp(79538) := x"0820";
    tmp(79539) := x"0000";
    tmp(79540) := x"0000";
    tmp(79541) := x"0000";
    tmp(79542) := x"0000";
    tmp(79543) := x"0000";
    tmp(79544) := x"0000";
    tmp(79545) := x"0000";
    tmp(79546) := x"0000";
    tmp(79547) := x"0000";
    tmp(79548) := x"0000";
    tmp(79549) := x"0000";
    tmp(79550) := x"0000";
    tmp(79551) := x"0000";
    tmp(79552) := x"0000";
    tmp(79553) := x"0000";
    tmp(79554) := x"0000";
    tmp(79555) := x"0000";
    tmp(79556) := x"0000";
    tmp(79557) := x"0000";
    tmp(79558) := x"0000";
    tmp(79559) := x"0000";
    tmp(79560) := x"0000";
    tmp(79561) := x"0000";
    tmp(79562) := x"0000";
    tmp(79563) := x"0000";
    tmp(79564) := x"0000";
    tmp(79565) := x"0000";
    tmp(79566) := x"0000";
    tmp(79567) := x"0000";
    tmp(79568) := x"0000";
    tmp(79569) := x"0000";
    tmp(79570) := x"0000";
    tmp(79571) := x"0000";
    tmp(79572) := x"0000";
    tmp(79573) := x"0000";
    tmp(79574) := x"0000";
    tmp(79575) := x"0000";
    tmp(79576) := x"0000";
    tmp(79577) := x"0000";
    tmp(79578) := x"0000";
    tmp(79579) := x"0000";
    tmp(79580) := x"0000";
    tmp(79581) := x"0000";
    tmp(79582) := x"0000";
    tmp(79583) := x"0000";
    tmp(79584) := x"0000";
    tmp(79585) := x"0000";
    tmp(79586) := x"0000";
    tmp(79587) := x"0000";
    tmp(79588) := x"0000";
    tmp(79589) := x"0000";
    tmp(79590) := x"0000";
    tmp(79591) := x"0000";
    tmp(79592) := x"0000";
    tmp(79593) := x"0000";
    tmp(79594) := x"0000";
    tmp(79595) := x"0000";
    tmp(79596) := x"0000";
    tmp(79597) := x"0000";
    tmp(79598) := x"0000";
    tmp(79599) := x"0000";
    tmp(79600) := x"0000";
    tmp(79601) := x"0000";
    tmp(79602) := x"0000";
    tmp(79603) := x"0000";
    tmp(79604) := x"0000";
    tmp(79605) := x"0000";
    tmp(79606) := x"0000";
    tmp(79607) := x"0000";
    tmp(79608) := x"0000";
    tmp(79609) := x"0000";
    tmp(79610) := x"0000";
    tmp(79611) := x"0000";
    tmp(79612) := x"0000";
    tmp(79613) := x"0000";
    tmp(79614) := x"0000";
    tmp(79615) := x"0000";
    tmp(79616) := x"0000";
    tmp(79617) := x"0000";
    tmp(79618) := x"0000";
    tmp(79619) := x"0000";
    tmp(79620) := x"0000";
    tmp(79621) := x"0000";
    tmp(79622) := x"0000";
    tmp(79623) := x"0000";
    tmp(79624) := x"0000";
    tmp(79625) := x"0000";
    tmp(79626) := x"0000";
    tmp(79627) := x"0000";
    tmp(79628) := x"0000";
    tmp(79629) := x"0000";
    tmp(79630) := x"0000";
    tmp(79631) := x"0000";
    tmp(79632) := x"0000";
    tmp(79633) := x"0000";
    tmp(79634) := x"0000";
    tmp(79635) := x"0000";
    tmp(79636) := x"0000";
    tmp(79637) := x"0000";
    tmp(79638) := x"0000";
    tmp(79639) := x"0000";
    tmp(79640) := x"0000";
    tmp(79641) := x"0000";
    tmp(79642) := x"0000";
    tmp(79643) := x"0000";
    tmp(79644) := x"0000";
    tmp(79645) := x"0000";
    tmp(79646) := x"0000";
    tmp(79647) := x"0000";
    tmp(79648) := x"0000";
    tmp(79649) := x"0000";
    tmp(79650) := x"0000";
    tmp(79651) := x"0000";
    tmp(79652) := x"0000";
    tmp(79653) := x"0000";
    tmp(79654) := x"0000";
    tmp(79655) := x"0000";
    tmp(79656) := x"0000";
    tmp(79657) := x"0000";
    tmp(79658) := x"0000";
    tmp(79659) := x"0000";
    tmp(79660) := x"0000";
    tmp(79661) := x"0000";
    tmp(79662) := x"0000";
    tmp(79663) := x"0000";
    tmp(79664) := x"0000";
    tmp(79665) := x"0000";
    tmp(79666) := x"0000";
    tmp(79667) := x"0000";
    tmp(79668) := x"0000";
    tmp(79669) := x"0000";
    tmp(79670) := x"0000";
    tmp(79671) := x"0000";
    tmp(79672) := x"0000";
    tmp(79673) := x"0000";
    tmp(79674) := x"0000";
    tmp(79675) := x"0000";
    tmp(79676) := x"0000";
    tmp(79677) := x"0000";
    tmp(79678) := x"0000";
    tmp(79679) := x"0000";
    tmp(79680) := x"0000";
    tmp(79681) := x"0020";
    tmp(79682) := x"0020";
    tmp(79683) := x"0020";
    tmp(79684) := x"0020";
    tmp(79685) := x"0020";
    tmp(79686) := x"0020";
    tmp(79687) := x"0020";
    tmp(79688) := x"0020";
    tmp(79689) := x"0020";
    tmp(79690) := x"0020";
    tmp(79691) := x"0020";
    tmp(79692) := x"0020";
    tmp(79693) := x"0020";
    tmp(79694) := x"0020";
    tmp(79695) := x"0020";
    tmp(79696) := x"0020";
    tmp(79697) := x"0020";
    tmp(79698) := x"0020";
    tmp(79699) := x"0020";
    tmp(79700) := x"0020";
    tmp(79701) := x"0020";
    tmp(79702) := x"0020";
    tmp(79703) := x"0020";
    tmp(79704) := x"0020";
    tmp(79705) := x"0020";
    tmp(79706) := x"0020";
    tmp(79707) := x"0020";
    tmp(79708) := x"0020";
    tmp(79709) := x"0020";
    tmp(79710) := x"0020";
    tmp(79711) := x"0020";
    tmp(79712) := x"0020";
    tmp(79713) := x"0020";
    tmp(79714) := x"0020";
    tmp(79715) := x"0820";
    tmp(79716) := x"0820";
    tmp(79717) := x"0820";
    tmp(79718) := x"0820";
    tmp(79719) := x"0820";
    tmp(79720) := x"0820";
    tmp(79721) := x"0820";
    tmp(79722) := x"0820";
    tmp(79723) := x"0820";
    tmp(79724) := x"0820";
    tmp(79725) := x"0820";
    tmp(79726) := x"0800";
    tmp(79727) := x"0800";
    tmp(79728) := x"0800";
    tmp(79729) := x"0800";
    tmp(79730) := x"0800";
    tmp(79731) := x"0800";
    tmp(79732) := x"0800";
    tmp(79733) := x"0800";
    tmp(79734) := x"1000";
    tmp(79735) := x"1000";
    tmp(79736) := x"1000";
    tmp(79737) := x"0800";
    tmp(79738) := x"0800";
    tmp(79739) := x"0800";
    tmp(79740) := x"1000";
    tmp(79741) := x"1000";
    tmp(79742) := x"1800";
    tmp(79743) := x"1000";
    tmp(79744) := x"1000";
    tmp(79745) := x"1000";
    tmp(79746) := x"1800";
    tmp(79747) := x"1800";
    tmp(79748) := x"1800";
    tmp(79749) := x"1800";
    tmp(79750) := x"1000";
    tmp(79751) := x"1000";
    tmp(79752) := x"1820";
    tmp(79753) := x"1820";
    tmp(79754) := x"1820";
    tmp(79755) := x"1020";
    tmp(79756) := x"0800";
    tmp(79757) := x"0000";
    tmp(79758) := x"0000";
    tmp(79759) := x"0000";
    tmp(79760) := x"0000";
    tmp(79761) := x"0000";
    tmp(79762) := x"0000";
    tmp(79763) := x"0000";
    tmp(79764) := x"0800";
    tmp(79765) := x"0800";
    tmp(79766) := x"0800";
    tmp(79767) := x"0800";
    tmp(79768) := x"0800";
    tmp(79769) := x"0800";
    tmp(79770) := x"0800";
    tmp(79771) := x"0800";
    tmp(79772) := x"0800";
    tmp(79773) := x"1000";
    tmp(79774) := x"0800";
    tmp(79775) := x"1000";
    tmp(79776) := x"1020";
    tmp(79777) := x"0820";
    tmp(79778) := x"0000";
    tmp(79779) := x"0000";
    tmp(79780) := x"0000";
    tmp(79781) := x"0000";
    tmp(79782) := x"0000";
    tmp(79783) := x"0000";
    tmp(79784) := x"0000";
    tmp(79785) := x"0000";
    tmp(79786) := x"0000";
    tmp(79787) := x"0000";
    tmp(79788) := x"0000";
    tmp(79789) := x"0000";
    tmp(79790) := x"0000";
    tmp(79791) := x"0000";
    tmp(79792) := x"0000";
    tmp(79793) := x"0000";
    tmp(79794) := x"0000";
    tmp(79795) := x"0000";
    tmp(79796) := x"0000";
    tmp(79797) := x"0000";
    tmp(79798) := x"0000";
    tmp(79799) := x"0000";
    tmp(79800) := x"0000";
    tmp(79801) := x"0000";
    tmp(79802) := x"0000";
    tmp(79803) := x"0000";
    tmp(79804) := x"0000";
    tmp(79805) := x"0000";
    tmp(79806) := x"0000";
    tmp(79807) := x"0000";
    tmp(79808) := x"0000";
    tmp(79809) := x"0000";
    tmp(79810) := x"0000";
    tmp(79811) := x"0000";
    tmp(79812) := x"0000";
    tmp(79813) := x"0000";
    tmp(79814) := x"0000";
    tmp(79815) := x"0000";
    tmp(79816) := x"0000";
    tmp(79817) := x"0000";
    tmp(79818) := x"0000";
    tmp(79819) := x"0000";
    tmp(79820) := x"0000";
    tmp(79821) := x"0000";
    tmp(79822) := x"0000";
    tmp(79823) := x"0000";
    tmp(79824) := x"0000";
    tmp(79825) := x"0000";
    tmp(79826) := x"0000";
    tmp(79827) := x"0000";
    tmp(79828) := x"0000";
    tmp(79829) := x"0000";
    tmp(79830) := x"0000";
    tmp(79831) := x"0000";
    tmp(79832) := x"0000";
    tmp(79833) := x"0000";
    tmp(79834) := x"0000";
    tmp(79835) := x"0000";
    tmp(79836) := x"0000";
    tmp(79837) := x"0000";
    tmp(79838) := x"0000";
    tmp(79839) := x"0000";
    tmp(79840) := x"0000";
    tmp(79841) := x"0000";
    tmp(79842) := x"0000";
    tmp(79843) := x"0000";
    tmp(79844) := x"0000";
    tmp(79845) := x"0000";
    tmp(79846) := x"0000";
    tmp(79847) := x"0000";
    tmp(79848) := x"0000";
    tmp(79849) := x"0000";
    tmp(79850) := x"0000";
    tmp(79851) := x"0000";
    tmp(79852) := x"0000";
    tmp(79853) := x"0000";
    tmp(79854) := x"0000";
    tmp(79855) := x"0000";
    tmp(79856) := x"0000";
    tmp(79857) := x"0000";
    tmp(79858) := x"0000";
    tmp(79859) := x"0000";
    tmp(79860) := x"0000";
    tmp(79861) := x"0000";
    tmp(79862) := x"0000";
    tmp(79863) := x"0000";
    tmp(79864) := x"0000";
    tmp(79865) := x"0000";
    tmp(79866) := x"0000";
    tmp(79867) := x"0000";
    tmp(79868) := x"0000";
    tmp(79869) := x"0000";
    tmp(79870) := x"0000";
    tmp(79871) := x"0000";
    tmp(79872) := x"0000";
    tmp(79873) := x"0000";
    tmp(79874) := x"0000";
    tmp(79875) := x"0000";
    tmp(79876) := x"0000";
    tmp(79877) := x"0000";
    tmp(79878) := x"0000";
    tmp(79879) := x"0000";
    tmp(79880) := x"0000";
    tmp(79881) := x"0000";
    tmp(79882) := x"0000";
    tmp(79883) := x"0000";
    tmp(79884) := x"0000";
    tmp(79885) := x"0000";
    tmp(79886) := x"0000";
    tmp(79887) := x"0000";
    tmp(79888) := x"0000";
    tmp(79889) := x"0000";
    tmp(79890) := x"0000";
    tmp(79891) := x"0000";
    tmp(79892) := x"0000";
    tmp(79893) := x"0000";
    tmp(79894) := x"0000";
    tmp(79895) := x"0000";
    tmp(79896) := x"0000";
    tmp(79897) := x"0000";
    tmp(79898) := x"0000";
    tmp(79899) := x"0000";
    tmp(79900) := x"0000";
    tmp(79901) := x"0000";
    tmp(79902) := x"0000";
    tmp(79903) := x"0000";
    tmp(79904) := x"0000";
    tmp(79905) := x"0000";
    tmp(79906) := x"0000";
    tmp(79907) := x"0000";
    tmp(79908) := x"0000";
    tmp(79909) := x"0000";
    tmp(79910) := x"0000";
    tmp(79911) := x"0000";
    tmp(79912) := x"0000";
    tmp(79913) := x"0000";
    tmp(79914) := x"0000";
    tmp(79915) := x"0000";
    tmp(79916) := x"0000";
    tmp(79917) := x"0000";
    tmp(79918) := x"0000";
    tmp(79919) := x"0000";
    tmp(79920) := x"0000";
    tmp(79921) := x"0020";
    tmp(79922) := x"0020";
    tmp(79923) := x"0020";
    tmp(79924) := x"0020";
    tmp(79925) := x"0020";
    tmp(79926) := x"0020";
    tmp(79927) := x"0020";
    tmp(79928) := x"0020";
    tmp(79929) := x"0020";
    tmp(79930) := x"0020";
    tmp(79931) := x"0020";
    tmp(79932) := x"0020";
    tmp(79933) := x"0020";
    tmp(79934) := x"0020";
    tmp(79935) := x"0020";
    tmp(79936) := x"0020";
    tmp(79937) := x"0020";
    tmp(79938) := x"0020";
    tmp(79939) := x"0020";
    tmp(79940) := x"0020";
    tmp(79941) := x"0020";
    tmp(79942) := x"0020";
    tmp(79943) := x"0020";
    tmp(79944) := x"0020";
    tmp(79945) := x"0020";
    tmp(79946) := x"0020";
    tmp(79947) := x"0020";
    tmp(79948) := x"0020";
    tmp(79949) := x"0020";
    tmp(79950) := x"0040";
    tmp(79951) := x"0040";
    tmp(79952) := x"0020";
    tmp(79953) := x"0020";
    tmp(79954) := x"0020";
    tmp(79955) := x"0020";
    tmp(79956) := x"0820";
    tmp(79957) := x"0820";
    tmp(79958) := x"0820";
    tmp(79959) := x"0820";
    tmp(79960) := x"0820";
    tmp(79961) := x"0820";
    tmp(79962) := x"0820";
    tmp(79963) := x"0820";
    tmp(79964) := x"0800";
    tmp(79965) := x"0800";
    tmp(79966) := x"0800";
    tmp(79967) := x"0800";
    tmp(79968) := x"0800";
    tmp(79969) := x"0800";
    tmp(79970) := x"0800";
    tmp(79971) := x"0800";
    tmp(79972) := x"0800";
    tmp(79973) := x"0800";
    tmp(79974) := x"1000";
    tmp(79975) := x"1000";
    tmp(79976) := x"1000";
    tmp(79977) := x"1000";
    tmp(79978) := x"0800";
    tmp(79979) := x"1000";
    tmp(79980) := x"1000";
    tmp(79981) := x"1000";
    tmp(79982) := x"1000";
    tmp(79983) := x"1000";
    tmp(79984) := x"1000";
    tmp(79985) := x"1000";
    tmp(79986) := x"1000";
    tmp(79987) := x"1000";
    tmp(79988) := x"1000";
    tmp(79989) := x"1800";
    tmp(79990) := x"1000";
    tmp(79991) := x"1000";
    tmp(79992) := x"1000";
    tmp(79993) := x"0800";
    tmp(79994) := x"0000";
    tmp(79995) := x"0000";
    tmp(79996) := x"0000";
    tmp(79997) := x"0000";
    tmp(79998) := x"0000";
    tmp(79999) := x"0000";
    tmp(80000) := x"0000";
    tmp(80001) := x"0000";
    tmp(80002) := x"0000";
    tmp(80003) := x"0800";
    tmp(80004) := x"1000";
    tmp(80005) := x"0800";
    tmp(80006) := x"0800";
    tmp(80007) := x"0800";
    tmp(80008) := x"0800";
    tmp(80009) := x"0800";
    tmp(80010) := x"0800";
    tmp(80011) := x"0800";
    tmp(80012) := x"1000";
    tmp(80013) := x"0800";
    tmp(80014) := x"0800";
    tmp(80015) := x"1020";
    tmp(80016) := x"0820";
    tmp(80017) := x"0000";
    tmp(80018) := x"0000";
    tmp(80019) := x"0000";
    tmp(80020) := x"0000";
    tmp(80021) := x"0000";
    tmp(80022) := x"0000";
    tmp(80023) := x"0000";
    tmp(80024) := x"0000";
    tmp(80025) := x"0000";
    tmp(80026) := x"0000";
    tmp(80027) := x"0000";
    tmp(80028) := x"0000";
    tmp(80029) := x"0000";
    tmp(80030) := x"0000";
    tmp(80031) := x"0000";
    tmp(80032) := x"0000";
    tmp(80033) := x"0000";
    tmp(80034) := x"0000";
    tmp(80035) := x"0000";
    tmp(80036) := x"0000";
    tmp(80037) := x"0000";
    tmp(80038) := x"0000";
    tmp(80039) := x"0000";
    tmp(80040) := x"0000";
    tmp(80041) := x"0000";
    tmp(80042) := x"0000";
    tmp(80043) := x"0000";
    tmp(80044) := x"0000";
    tmp(80045) := x"0000";
    tmp(80046) := x"0000";
    tmp(80047) := x"0000";
    tmp(80048) := x"0000";
    tmp(80049) := x"0000";
    tmp(80050) := x"0000";
    tmp(80051) := x"0000";
    tmp(80052) := x"0000";
    tmp(80053) := x"0000";
    tmp(80054) := x"0000";
    tmp(80055) := x"0000";
    tmp(80056) := x"0000";
    tmp(80057) := x"0000";
    tmp(80058) := x"0000";
    tmp(80059) := x"0000";
    tmp(80060) := x"0000";
    tmp(80061) := x"0000";
    tmp(80062) := x"0000";
    tmp(80063) := x"0000";
    tmp(80064) := x"0000";
    tmp(80065) := x"0000";
    tmp(80066) := x"0000";
    tmp(80067) := x"0000";
    tmp(80068) := x"0000";
    tmp(80069) := x"0000";
    tmp(80070) := x"0000";
    tmp(80071) := x"0000";
    tmp(80072) := x"0000";
    tmp(80073) := x"0000";
    tmp(80074) := x"0000";
    tmp(80075) := x"0000";
    tmp(80076) := x"0000";
    tmp(80077) := x"0000";
    tmp(80078) := x"0000";
    tmp(80079) := x"0000";
    tmp(80080) := x"0000";
    tmp(80081) := x"0000";
    tmp(80082) := x"0000";
    tmp(80083) := x"0000";
    tmp(80084) := x"0000";
    tmp(80085) := x"0000";
    tmp(80086) := x"0000";
    tmp(80087) := x"0000";
    tmp(80088) := x"0000";
    tmp(80089) := x"0000";
    tmp(80090) := x"0000";
    tmp(80091) := x"0000";
    tmp(80092) := x"0000";
    tmp(80093) := x"0000";
    tmp(80094) := x"0000";
    tmp(80095) := x"0000";
    tmp(80096) := x"0000";
    tmp(80097) := x"0000";
    tmp(80098) := x"0000";
    tmp(80099) := x"0000";
    tmp(80100) := x"0000";
    tmp(80101) := x"0000";
    tmp(80102) := x"0000";
    tmp(80103) := x"0000";
    tmp(80104) := x"0000";
    tmp(80105) := x"0000";
    tmp(80106) := x"0000";
    tmp(80107) := x"0000";
    tmp(80108) := x"0000";
    tmp(80109) := x"0000";
    tmp(80110) := x"0000";
    tmp(80111) := x"0000";
    tmp(80112) := x"0000";
    tmp(80113) := x"0000";
    tmp(80114) := x"0000";
    tmp(80115) := x"0000";
    tmp(80116) := x"0000";
    tmp(80117) := x"0000";
    tmp(80118) := x"0000";
    tmp(80119) := x"0000";
    tmp(80120) := x"0000";
    tmp(80121) := x"0000";
    tmp(80122) := x"0000";
    tmp(80123) := x"0000";
    tmp(80124) := x"0000";
    tmp(80125) := x"0000";
    tmp(80126) := x"0000";
    tmp(80127) := x"0000";
    tmp(80128) := x"0000";
    tmp(80129) := x"0000";
    tmp(80130) := x"0000";
    tmp(80131) := x"0000";
    tmp(80132) := x"0000";
    tmp(80133) := x"0000";
    tmp(80134) := x"0000";
    tmp(80135) := x"0000";
    tmp(80136) := x"0000";
    tmp(80137) := x"0000";
    tmp(80138) := x"0000";
    tmp(80139) := x"0000";
    tmp(80140) := x"0000";
    tmp(80141) := x"0000";
    tmp(80142) := x"0000";
    tmp(80143) := x"0000";
    tmp(80144) := x"0000";
    tmp(80145) := x"0000";
    tmp(80146) := x"0000";
    tmp(80147) := x"0000";
    tmp(80148) := x"0000";
    tmp(80149) := x"0000";
    tmp(80150) := x"0000";
    tmp(80151) := x"0000";
    tmp(80152) := x"0000";
    tmp(80153) := x"0000";
    tmp(80154) := x"0000";
    tmp(80155) := x"0000";
    tmp(80156) := x"0000";
    tmp(80157) := x"0000";
    tmp(80158) := x"0000";
    tmp(80159) := x"0000";
    tmp(80160) := x"0000";
    tmp(80161) := x"0020";
    tmp(80162) := x"0020";
    tmp(80163) := x"0020";
    tmp(80164) := x"0020";
    tmp(80165) := x"0020";
    tmp(80166) := x"0020";
    tmp(80167) := x"0020";
    tmp(80168) := x"0020";
    tmp(80169) := x"0020";
    tmp(80170) := x"0020";
    tmp(80171) := x"0020";
    tmp(80172) := x"0020";
    tmp(80173) := x"0020";
    tmp(80174) := x"0020";
    tmp(80175) := x"0020";
    tmp(80176) := x"0020";
    tmp(80177) := x"0020";
    tmp(80178) := x"0020";
    tmp(80179) := x"0020";
    tmp(80180) := x"0020";
    tmp(80181) := x"0020";
    tmp(80182) := x"0020";
    tmp(80183) := x"0020";
    tmp(80184) := x"0020";
    tmp(80185) := x"0020";
    tmp(80186) := x"0020";
    tmp(80187) := x"0020";
    tmp(80188) := x"0020";
    tmp(80189) := x"0020";
    tmp(80190) := x"0020";
    tmp(80191) := x"0020";
    tmp(80192) := x"0020";
    tmp(80193) := x"0020";
    tmp(80194) := x"0020";
    tmp(80195) := x"0020";
    tmp(80196) := x"0820";
    tmp(80197) := x"0820";
    tmp(80198) := x"0820";
    tmp(80199) := x"0820";
    tmp(80200) := x"0820";
    tmp(80201) := x"0820";
    tmp(80202) := x"0800";
    tmp(80203) := x"0800";
    tmp(80204) := x"0800";
    tmp(80205) := x"0800";
    tmp(80206) := x"0800";
    tmp(80207) := x"0800";
    tmp(80208) := x"0800";
    tmp(80209) := x"0800";
    tmp(80210) := x"0800";
    tmp(80211) := x"0800";
    tmp(80212) := x"0800";
    tmp(80213) := x"0800";
    tmp(80214) := x"0800";
    tmp(80215) := x"1000";
    tmp(80216) := x"1000";
    tmp(80217) := x"1000";
    tmp(80218) := x"0800";
    tmp(80219) := x"0800";
    tmp(80220) := x"0800";
    tmp(80221) := x"1000";
    tmp(80222) := x"1000";
    tmp(80223) := x"1000";
    tmp(80224) := x"1000";
    tmp(80225) := x"1000";
    tmp(80226) := x"1000";
    tmp(80227) := x"1000";
    tmp(80228) := x"1000";
    tmp(80229) := x"1000";
    tmp(80230) := x"0800";
    tmp(80231) := x"0800";
    tmp(80232) := x"0000";
    tmp(80233) := x"0000";
    tmp(80234) := x"0000";
    tmp(80235) := x"0000";
    tmp(80236) := x"0000";
    tmp(80237) := x"0000";
    tmp(80238) := x"0000";
    tmp(80239) := x"0000";
    tmp(80240) := x"0000";
    tmp(80241) := x"0000";
    tmp(80242) := x"0800";
    tmp(80243) := x"0800";
    tmp(80244) := x"0800";
    tmp(80245) := x"0000";
    tmp(80246) := x"0800";
    tmp(80247) := x"0800";
    tmp(80248) := x"1000";
    tmp(80249) := x"0800";
    tmp(80250) := x"0800";
    tmp(80251) := x"1000";
    tmp(80252) := x"1000";
    tmp(80253) := x"1000";
    tmp(80254) := x"1020";
    tmp(80255) := x"0820";
    tmp(80256) := x"0000";
    tmp(80257) := x"0000";
    tmp(80258) := x"0000";
    tmp(80259) := x"0000";
    tmp(80260) := x"0000";
    tmp(80261) := x"0000";
    tmp(80262) := x"0000";
    tmp(80263) := x"0000";
    tmp(80264) := x"0000";
    tmp(80265) := x"0000";
    tmp(80266) := x"0000";
    tmp(80267) := x"0000";
    tmp(80268) := x"0000";
    tmp(80269) := x"0000";
    tmp(80270) := x"0000";
    tmp(80271) := x"0000";
    tmp(80272) := x"0000";
    tmp(80273) := x"0000";
    tmp(80274) := x"0000";
    tmp(80275) := x"0000";
    tmp(80276) := x"0000";
    tmp(80277) := x"0000";
    tmp(80278) := x"0000";
    tmp(80279) := x"0000";
    tmp(80280) := x"0000";
    tmp(80281) := x"0000";
    tmp(80282) := x"0000";
    tmp(80283) := x"0000";
    tmp(80284) := x"0000";
    tmp(80285) := x"0000";
    tmp(80286) := x"0000";
    tmp(80287) := x"0000";
    tmp(80288) := x"0000";
    tmp(80289) := x"0000";
    tmp(80290) := x"0000";
    tmp(80291) := x"0000";
    tmp(80292) := x"0000";
    tmp(80293) := x"0000";
    tmp(80294) := x"0000";
    tmp(80295) := x"0000";
    tmp(80296) := x"0000";
    tmp(80297) := x"0000";
    tmp(80298) := x"0000";
    tmp(80299) := x"0000";
    tmp(80300) := x"0000";
    tmp(80301) := x"0000";
    tmp(80302) := x"0000";
    tmp(80303) := x"0000";
    tmp(80304) := x"0000";
    tmp(80305) := x"0000";
    tmp(80306) := x"0000";
    tmp(80307) := x"0000";
    tmp(80308) := x"0000";
    tmp(80309) := x"0000";
    tmp(80310) := x"0000";
    tmp(80311) := x"0000";
    tmp(80312) := x"0000";
    tmp(80313) := x"0000";
    tmp(80314) := x"0000";
    tmp(80315) := x"0000";
    tmp(80316) := x"0000";
    tmp(80317) := x"0000";
    tmp(80318) := x"0000";
    tmp(80319) := x"0000";
    tmp(80320) := x"0000";
    tmp(80321) := x"0000";
    tmp(80322) := x"0000";
    tmp(80323) := x"0000";
    tmp(80324) := x"0000";
    tmp(80325) := x"0000";
    tmp(80326) := x"0000";
    tmp(80327) := x"0000";
    tmp(80328) := x"0000";
    tmp(80329) := x"0000";
    tmp(80330) := x"0000";
    tmp(80331) := x"0000";
    tmp(80332) := x"0000";
    tmp(80333) := x"0000";
    tmp(80334) := x"0000";
    tmp(80335) := x"0000";
    tmp(80336) := x"0000";
    tmp(80337) := x"0000";
    tmp(80338) := x"0000";
    tmp(80339) := x"0000";
    tmp(80340) := x"0000";
    tmp(80341) := x"0000";
    tmp(80342) := x"0000";
    tmp(80343) := x"0000";
    tmp(80344) := x"0000";
    tmp(80345) := x"0000";
    tmp(80346) := x"0000";
    tmp(80347) := x"0000";
    tmp(80348) := x"0000";
    tmp(80349) := x"0000";
    tmp(80350) := x"0000";
    tmp(80351) := x"0000";
    tmp(80352) := x"0000";
    tmp(80353) := x"0000";
    tmp(80354) := x"0000";
    tmp(80355) := x"0000";
    tmp(80356) := x"0000";
    tmp(80357) := x"0000";
    tmp(80358) := x"0000";
    tmp(80359) := x"0000";
    tmp(80360) := x"0000";
    tmp(80361) := x"0000";
    tmp(80362) := x"0000";
    tmp(80363) := x"0000";
    tmp(80364) := x"0000";
    tmp(80365) := x"0000";
    tmp(80366) := x"0000";
    tmp(80367) := x"0000";
    tmp(80368) := x"0000";
    tmp(80369) := x"0000";
    tmp(80370) := x"0000";
    tmp(80371) := x"0000";
    tmp(80372) := x"0000";
    tmp(80373) := x"0000";
    tmp(80374) := x"0000";
    tmp(80375) := x"0000";
    tmp(80376) := x"0000";
    tmp(80377) := x"0000";
    tmp(80378) := x"0000";
    tmp(80379) := x"0000";
    tmp(80380) := x"0000";
    tmp(80381) := x"0000";
    tmp(80382) := x"0000";
    tmp(80383) := x"0000";
    tmp(80384) := x"0000";
    tmp(80385) := x"0000";
    tmp(80386) := x"0000";
    tmp(80387) := x"0000";
    tmp(80388) := x"0000";
    tmp(80389) := x"0000";
    tmp(80390) := x"0000";
    tmp(80391) := x"0000";
    tmp(80392) := x"0000";
    tmp(80393) := x"0000";
    tmp(80394) := x"0000";
    tmp(80395) := x"0000";
    tmp(80396) := x"0000";
    tmp(80397) := x"0000";
    tmp(80398) := x"0000";
    tmp(80399) := x"0000";
    tmp(80400) := x"0000";
    tmp(80401) := x"0000";
    tmp(80402) := x"0000";
    tmp(80403) := x"0000";
    tmp(80404) := x"0000";
    tmp(80405) := x"0020";
    tmp(80406) := x"0020";
    tmp(80407) := x"0020";
    tmp(80408) := x"0020";
    tmp(80409) := x"0020";
    tmp(80410) := x"0020";
    tmp(80411) := x"0020";
    tmp(80412) := x"0020";
    tmp(80413) := x"0020";
    tmp(80414) := x"0020";
    tmp(80415) := x"0020";
    tmp(80416) := x"0020";
    tmp(80417) := x"0020";
    tmp(80418) := x"0020";
    tmp(80419) := x"0020";
    tmp(80420) := x"0020";
    tmp(80421) := x"0020";
    tmp(80422) := x"0020";
    tmp(80423) := x"0020";
    tmp(80424) := x"0020";
    tmp(80425) := x"0020";
    tmp(80426) := x"0020";
    tmp(80427) := x"0020";
    tmp(80428) := x"0020";
    tmp(80429) := x"0020";
    tmp(80430) := x"0020";
    tmp(80431) := x"0000";
    tmp(80432) := x"0000";
    tmp(80433) := x"0000";
    tmp(80434) := x"0000";
    tmp(80435) := x"0020";
    tmp(80436) := x"0800";
    tmp(80437) := x"0800";
    tmp(80438) := x"0800";
    tmp(80439) := x"0800";
    tmp(80440) := x"0000";
    tmp(80441) := x"0000";
    tmp(80442) := x"0000";
    tmp(80443) := x"0800";
    tmp(80444) := x"0800";
    tmp(80445) := x"0800";
    tmp(80446) := x"0800";
    tmp(80447) := x"0800";
    tmp(80448) := x"0800";
    tmp(80449) := x"0800";
    tmp(80450) := x"0800";
    tmp(80451) := x"0800";
    tmp(80452) := x"0800";
    tmp(80453) := x"0800";
    tmp(80454) := x"0800";
    tmp(80455) := x"0800";
    tmp(80456) := x"0800";
    tmp(80457) := x"0800";
    tmp(80458) := x"0800";
    tmp(80459) := x"0800";
    tmp(80460) := x"0800";
    tmp(80461) := x"0800";
    tmp(80462) := x"1000";
    tmp(80463) := x"1000";
    tmp(80464) := x"1000";
    tmp(80465) := x"1000";
    tmp(80466) := x"1000";
    tmp(80467) := x"1000";
    tmp(80468) := x"0800";
    tmp(80469) := x"0800";
    tmp(80470) := x"0000";
    tmp(80471) := x"0000";
    tmp(80472) := x"0000";
    tmp(80473) := x"0000";
    tmp(80474) := x"0000";
    tmp(80475) := x"0000";
    tmp(80476) := x"0800";
    tmp(80477) := x"0000";
    tmp(80478) := x"0000";
    tmp(80479) := x"0800";
    tmp(80480) := x"0800";
    tmp(80481) := x"0800";
    tmp(80482) := x"0800";
    tmp(80483) := x"0000";
    tmp(80484) := x"0800";
    tmp(80485) := x"0800";
    tmp(80486) := x"0800";
    tmp(80487) := x"0800";
    tmp(80488) := x"0800";
    tmp(80489) := x"1000";
    tmp(80490) := x"1000";
    tmp(80491) := x"1000";
    tmp(80492) := x"1000";
    tmp(80493) := x"1020";
    tmp(80494) := x"0820";
    tmp(80495) := x"0000";
    tmp(80496) := x"0000";
    tmp(80497) := x"0000";
    tmp(80498) := x"0000";
    tmp(80499) := x"0000";
    tmp(80500) := x"0000";
    tmp(80501) := x"0000";
    tmp(80502) := x"0000";
    tmp(80503) := x"0000";
    tmp(80504) := x"0000";
    tmp(80505) := x"0000";
    tmp(80506) := x"0000";
    tmp(80507) := x"0000";
    tmp(80508) := x"0000";
    tmp(80509) := x"0000";
    tmp(80510) := x"0000";
    tmp(80511) := x"0000";
    tmp(80512) := x"0000";
    tmp(80513) := x"0000";
    tmp(80514) := x"0000";
    tmp(80515) := x"0000";
    tmp(80516) := x"0000";
    tmp(80517) := x"0000";
    tmp(80518) := x"0000";
    tmp(80519) := x"0000";
    tmp(80520) := x"0000";
    tmp(80521) := x"0000";
    tmp(80522) := x"0000";
    tmp(80523) := x"0000";
    tmp(80524) := x"0000";
    tmp(80525) := x"0000";
    tmp(80526) := x"0000";
    tmp(80527) := x"0000";
    tmp(80528) := x"0000";
    tmp(80529) := x"0000";
    tmp(80530) := x"0000";
    tmp(80531) := x"0000";
    tmp(80532) := x"0000";
    tmp(80533) := x"0000";
    tmp(80534) := x"0000";
    tmp(80535) := x"0000";
    tmp(80536) := x"0000";
    tmp(80537) := x"0000";
    tmp(80538) := x"0000";
    tmp(80539) := x"0000";
    tmp(80540) := x"0000";
    tmp(80541) := x"0000";
    tmp(80542) := x"0000";
    tmp(80543) := x"0000";
    tmp(80544) := x"0000";
    tmp(80545) := x"0000";
    tmp(80546) := x"0000";
    tmp(80547) := x"0000";
    tmp(80548) := x"0000";
    tmp(80549) := x"0000";
    tmp(80550) := x"0000";
    tmp(80551) := x"0000";
    tmp(80552) := x"0000";
    tmp(80553) := x"0000";
    tmp(80554) := x"0000";
    tmp(80555) := x"0000";
    tmp(80556) := x"0000";
    tmp(80557) := x"0000";
    tmp(80558) := x"0000";
    tmp(80559) := x"0000";
    tmp(80560) := x"0000";
    tmp(80561) := x"0000";
    tmp(80562) := x"0000";
    tmp(80563) := x"0000";
    tmp(80564) := x"0000";
    tmp(80565) := x"0000";
    tmp(80566) := x"0000";
    tmp(80567) := x"0000";
    tmp(80568) := x"0000";
    tmp(80569) := x"0000";
    tmp(80570) := x"0000";
    tmp(80571) := x"0000";
    tmp(80572) := x"0000";
    tmp(80573) := x"0000";
    tmp(80574) := x"0000";
    tmp(80575) := x"0000";
    tmp(80576) := x"0000";
    tmp(80577) := x"0000";
    tmp(80578) := x"0000";
    tmp(80579) := x"0000";
    tmp(80580) := x"0000";
    tmp(80581) := x"0000";
    tmp(80582) := x"0000";
    tmp(80583) := x"0000";
    tmp(80584) := x"0000";
    tmp(80585) := x"0000";
    tmp(80586) := x"0000";
    tmp(80587) := x"0000";
    tmp(80588) := x"0000";
    tmp(80589) := x"0000";
    tmp(80590) := x"0000";
    tmp(80591) := x"0000";
    tmp(80592) := x"0000";
    tmp(80593) := x"0000";
    tmp(80594) := x"0000";
    tmp(80595) := x"0000";
    tmp(80596) := x"0000";
    tmp(80597) := x"0000";
    tmp(80598) := x"0000";
    tmp(80599) := x"0000";
    tmp(80600) := x"0000";
    tmp(80601) := x"0000";
    tmp(80602) := x"0000";
    tmp(80603) := x"0000";
    tmp(80604) := x"0000";
    tmp(80605) := x"0000";
    tmp(80606) := x"0000";
    tmp(80607) := x"0000";
    tmp(80608) := x"0000";
    tmp(80609) := x"0000";
    tmp(80610) := x"0000";
    tmp(80611) := x"0000";
    tmp(80612) := x"0000";
    tmp(80613) := x"0000";
    tmp(80614) := x"0000";
    tmp(80615) := x"0000";
    tmp(80616) := x"0000";
    tmp(80617) := x"0000";
    tmp(80618) := x"0000";
    tmp(80619) := x"0000";
    tmp(80620) := x"0000";
    tmp(80621) := x"0000";
    tmp(80622) := x"0000";
    tmp(80623) := x"0000";
    tmp(80624) := x"0000";
    tmp(80625) := x"0000";
    tmp(80626) := x"0000";
    tmp(80627) := x"0000";
    tmp(80628) := x"0000";
    tmp(80629) := x"0000";
    tmp(80630) := x"0000";
    tmp(80631) := x"0000";
    tmp(80632) := x"0000";
    tmp(80633) := x"0000";
    tmp(80634) := x"0000";
    tmp(80635) := x"0000";
    tmp(80636) := x"0000";
    tmp(80637) := x"0000";
    tmp(80638) := x"0000";
    tmp(80639) := x"0000";
    tmp(80640) := x"0000";
    tmp(80641) := x"0000";
    tmp(80642) := x"0000";
    tmp(80643) := x"0000";
    tmp(80644) := x"0000";
    tmp(80645) := x"0000";
    tmp(80646) := x"0000";
    tmp(80647) := x"0000";
    tmp(80648) := x"0000";
    tmp(80649) := x"0000";
    tmp(80650) := x"0000";
    tmp(80651) := x"0000";
    tmp(80652) := x"0000";
    tmp(80653) := x"0000";
    tmp(80654) := x"0000";
    tmp(80655) := x"0000";
    tmp(80656) := x"0000";
    tmp(80657) := x"0000";
    tmp(80658) := x"0000";
    tmp(80659) := x"0000";
    tmp(80660) := x"0000";
    tmp(80661) := x"0000";
    tmp(80662) := x"0000";
    tmp(80663) := x"0020";
    tmp(80664) := x"0020";
    tmp(80665) := x"0020";
    tmp(80666) := x"0020";
    tmp(80667) := x"0020";
    tmp(80668) := x"0020";
    tmp(80669) := x"0000";
    tmp(80670) := x"0800";
    tmp(80671) := x"0000";
    tmp(80672) := x"0000";
    tmp(80673) := x"0000";
    tmp(80674) := x"0020";
    tmp(80675) := x"0820";
    tmp(80676) := x"0800";
    tmp(80677) := x"0800";
    tmp(80678) := x"0800";
    tmp(80679) := x"0800";
    tmp(80680) := x"0000";
    tmp(80681) := x"0000";
    tmp(80682) := x"0800";
    tmp(80683) := x"0800";
    tmp(80684) := x"0800";
    tmp(80685) := x"0800";
    tmp(80686) := x"0800";
    tmp(80687) := x"0800";
    tmp(80688) := x"0800";
    tmp(80689) := x"0800";
    tmp(80690) := x"0800";
    tmp(80691) := x"0800";
    tmp(80692) := x"0800";
    tmp(80693) := x"0800";
    tmp(80694) := x"0800";
    tmp(80695) := x"0800";
    tmp(80696) := x"0800";
    tmp(80697) := x"0800";
    tmp(80698) := x"1000";
    tmp(80699) := x"1000";
    tmp(80700) := x"0800";
    tmp(80701) := x"0800";
    tmp(80702) := x"1000";
    tmp(80703) := x"1000";
    tmp(80704) := x"0800";
    tmp(80705) := x"0800";
    tmp(80706) := x"0800";
    tmp(80707) := x"0800";
    tmp(80708) := x"0800";
    tmp(80709) := x"0000";
    tmp(80710) := x"0000";
    tmp(80711) := x"0000";
    tmp(80712) := x"0000";
    tmp(80713) := x"0000";
    tmp(80714) := x"0800";
    tmp(80715) := x"0000";
    tmp(80716) := x"0000";
    tmp(80717) := x"0800";
    tmp(80718) := x"0800";
    tmp(80719) := x"0800";
    tmp(80720) := x"0000";
    tmp(80721) := x"0000";
    tmp(80722) := x"0000";
    tmp(80723) := x"0000";
    tmp(80724) := x"0000";
    tmp(80725) := x"0000";
    tmp(80726) := x"0800";
    tmp(80727) := x"0800";
    tmp(80728) := x"0800";
    tmp(80729) := x"1000";
    tmp(80730) := x"1000";
    tmp(80731) := x"1020";
    tmp(80732) := x"1020";
    tmp(80733) := x"0820";
    tmp(80734) := x"0000";
    tmp(80735) := x"0000";
    tmp(80736) := x"0000";
    tmp(80737) := x"0000";
    tmp(80738) := x"0000";
    tmp(80739) := x"0000";
    tmp(80740) := x"0000";
    tmp(80741) := x"0000";
    tmp(80742) := x"0000";
    tmp(80743) := x"0000";
    tmp(80744) := x"0000";
    tmp(80745) := x"0000";
    tmp(80746) := x"0000";
    tmp(80747) := x"0000";
    tmp(80748) := x"0000";
    tmp(80749) := x"0000";
    tmp(80750) := x"0000";
    tmp(80751) := x"0000";
    tmp(80752) := x"0000";
    tmp(80753) := x"0000";
    tmp(80754) := x"0000";
    tmp(80755) := x"0000";
    tmp(80756) := x"0000";
    tmp(80757) := x"0000";
    tmp(80758) := x"0000";
    tmp(80759) := x"0000";
    tmp(80760) := x"0000";
    tmp(80761) := x"0000";
    tmp(80762) := x"0000";
    tmp(80763) := x"0000";
    tmp(80764) := x"0000";
    tmp(80765) := x"0000";
    tmp(80766) := x"0000";
    tmp(80767) := x"0000";
    tmp(80768) := x"0000";
    tmp(80769) := x"0000";
    tmp(80770) := x"0000";
    tmp(80771) := x"0000";
    tmp(80772) := x"0000";
    tmp(80773) := x"0000";
    tmp(80774) := x"0000";
    tmp(80775) := x"0000";
    tmp(80776) := x"0000";
    tmp(80777) := x"0000";
    tmp(80778) := x"0000";
    tmp(80779) := x"0000";
    tmp(80780) := x"0000";
    tmp(80781) := x"0000";
    tmp(80782) := x"0000";
    tmp(80783) := x"0000";
    tmp(80784) := x"0000";
    tmp(80785) := x"0000";
    tmp(80786) := x"0000";
    tmp(80787) := x"0000";
    tmp(80788) := x"0000";
    tmp(80789) := x"0000";
    tmp(80790) := x"0000";
    tmp(80791) := x"0000";
    tmp(80792) := x"0000";
    tmp(80793) := x"0000";
    tmp(80794) := x"0000";
    tmp(80795) := x"0000";
    tmp(80796) := x"0000";
    tmp(80797) := x"0000";
    tmp(80798) := x"0000";
    tmp(80799) := x"0000";
    tmp(80800) := x"0000";
    tmp(80801) := x"0000";
    tmp(80802) := x"0000";
    tmp(80803) := x"0000";
    tmp(80804) := x"0000";
    tmp(80805) := x"0000";
    tmp(80806) := x"0000";
    tmp(80807) := x"0000";
    tmp(80808) := x"0000";
    tmp(80809) := x"0000";
    tmp(80810) := x"0000";
    tmp(80811) := x"0000";
    tmp(80812) := x"0000";
    tmp(80813) := x"0000";
    tmp(80814) := x"0000";
    tmp(80815) := x"0000";
    tmp(80816) := x"0000";
    tmp(80817) := x"0000";
    tmp(80818) := x"0000";
    tmp(80819) := x"0000";
    tmp(80820) := x"0000";
    tmp(80821) := x"0000";
    tmp(80822) := x"0000";
    tmp(80823) := x"0000";
    tmp(80824) := x"0000";
    tmp(80825) := x"0000";
    tmp(80826) := x"0000";
    tmp(80827) := x"0000";
    tmp(80828) := x"0000";
    tmp(80829) := x"0000";
    tmp(80830) := x"0000";
    tmp(80831) := x"0000";
    tmp(80832) := x"0000";
    tmp(80833) := x"0000";
    tmp(80834) := x"0000";
    tmp(80835) := x"0000";
    tmp(80836) := x"0000";
    tmp(80837) := x"0000";
    tmp(80838) := x"0000";
    tmp(80839) := x"0000";
    tmp(80840) := x"0000";
    tmp(80841) := x"0000";
    tmp(80842) := x"0000";
    tmp(80843) := x"0000";
    tmp(80844) := x"0000";
    tmp(80845) := x"0000";
    tmp(80846) := x"0000";
    tmp(80847) := x"0000";
    tmp(80848) := x"0000";
    tmp(80849) := x"0000";
    tmp(80850) := x"0000";
    tmp(80851) := x"0000";
    tmp(80852) := x"0000";
    tmp(80853) := x"0000";
    tmp(80854) := x"0000";
    tmp(80855) := x"0000";
    tmp(80856) := x"0000";
    tmp(80857) := x"0000";
    tmp(80858) := x"0000";
    tmp(80859) := x"0000";
    tmp(80860) := x"0000";
    tmp(80861) := x"0000";
    tmp(80862) := x"0000";
    tmp(80863) := x"0000";
    tmp(80864) := x"0000";
    tmp(80865) := x"0000";
    tmp(80866) := x"0000";
    tmp(80867) := x"0000";
    tmp(80868) := x"0000";
    tmp(80869) := x"0000";
    tmp(80870) := x"0000";
    tmp(80871) := x"0000";
    tmp(80872) := x"0000";
    tmp(80873) := x"0000";
    tmp(80874) := x"0000";
    tmp(80875) := x"0000";
    tmp(80876) := x"0000";
    tmp(80877) := x"0000";
    tmp(80878) := x"0000";
    tmp(80879) := x"0000";
    tmp(80880) := x"0000";
    tmp(80881) := x"0000";
    tmp(80882) := x"0000";
    tmp(80883) := x"0000";
    tmp(80884) := x"0000";
    tmp(80885) := x"0000";
    tmp(80886) := x"0000";
    tmp(80887) := x"0000";
    tmp(80888) := x"0000";
    tmp(80889) := x"0000";
    tmp(80890) := x"0000";
    tmp(80891) := x"0000";
    tmp(80892) := x"0000";
    tmp(80893) := x"0000";
    tmp(80894) := x"0000";
    tmp(80895) := x"0000";
    tmp(80896) := x"0000";
    tmp(80897) := x"0000";
    tmp(80898) := x"0000";
    tmp(80899) := x"0020";
    tmp(80900) := x"0020";
    tmp(80901) := x"0020";
    tmp(80902) := x"0020";
    tmp(80903) := x"0020";
    tmp(80904) := x"0020";
    tmp(80905) := x"0020";
    tmp(80906) := x"0020";
    tmp(80907) := x"0020";
    tmp(80908) := x"0020";
    tmp(80909) := x"0000";
    tmp(80910) := x"0800";
    tmp(80911) := x"0800";
    tmp(80912) := x"0800";
    tmp(80913) := x"0000";
    tmp(80914) := x"0000";
    tmp(80915) := x"0000";
    tmp(80916) := x"0000";
    tmp(80917) := x"0800";
    tmp(80918) := x"0800";
    tmp(80919) := x"0800";
    tmp(80920) := x"0800";
    tmp(80921) := x"0800";
    tmp(80922) := x"0800";
    tmp(80923) := x"0800";
    tmp(80924) := x"0800";
    tmp(80925) := x"0800";
    tmp(80926) := x"0800";
    tmp(80927) := x"0800";
    tmp(80928) := x"0800";
    tmp(80929) := x"0800";
    tmp(80930) := x"0800";
    tmp(80931) := x"0800";
    tmp(80932) := x"0800";
    tmp(80933) := x"0800";
    tmp(80934) := x"0800";
    tmp(80935) := x"1000";
    tmp(80936) := x"1000";
    tmp(80937) := x"1000";
    tmp(80938) := x"1000";
    tmp(80939) := x"0800";
    tmp(80940) := x"0800";
    tmp(80941) := x"0800";
    tmp(80942) := x"1000";
    tmp(80943) := x"1000";
    tmp(80944) := x"0800";
    tmp(80945) := x"0800";
    tmp(80946) := x"0800";
    tmp(80947) := x"0000";
    tmp(80948) := x"0000";
    tmp(80949) := x"0000";
    tmp(80950) := x"0000";
    tmp(80951) := x"0000";
    tmp(80952) := x"0800";
    tmp(80953) := x"0800";
    tmp(80954) := x"0000";
    tmp(80955) := x"0000";
    tmp(80956) := x"0800";
    tmp(80957) := x"0800";
    tmp(80958) := x"0000";
    tmp(80959) := x"0000";
    tmp(80960) := x"0000";
    tmp(80961) := x"0000";
    tmp(80962) := x"0000";
    tmp(80963) := x"0000";
    tmp(80964) := x"0000";
    tmp(80965) := x"0000";
    tmp(80966) := x"0000";
    tmp(80967) := x"0800";
    tmp(80968) := x"1000";
    tmp(80969) := x"1000";
    tmp(80970) := x"1020";
    tmp(80971) := x"0820";
    tmp(80972) := x"0000";
    tmp(80973) := x"0000";
    tmp(80974) := x"0000";
    tmp(80975) := x"0000";
    tmp(80976) := x"0000";
    tmp(80977) := x"0000";
    tmp(80978) := x"0000";
    tmp(80979) := x"0000";
    tmp(80980) := x"0000";
    tmp(80981) := x"0000";
    tmp(80982) := x"0000";
    tmp(80983) := x"0000";
    tmp(80984) := x"0000";
    tmp(80985) := x"0000";
    tmp(80986) := x"0000";
    tmp(80987) := x"0000";
    tmp(80988) := x"0000";
    tmp(80989) := x"0000";
    tmp(80990) := x"0000";
    tmp(80991) := x"0000";
    tmp(80992) := x"0000";
    tmp(80993) := x"0000";
    tmp(80994) := x"0000";
    tmp(80995) := x"0000";
    tmp(80996) := x"0000";
    tmp(80997) := x"0000";
    tmp(80998) := x"0000";
    tmp(80999) := x"0000";
    tmp(81000) := x"0000";
    tmp(81001) := x"0000";
    tmp(81002) := x"0000";
    tmp(81003) := x"0000";
    tmp(81004) := x"0000";
    tmp(81005) := x"0000";
    tmp(81006) := x"0000";
    tmp(81007) := x"0000";
    tmp(81008) := x"0000";
    tmp(81009) := x"0000";
    tmp(81010) := x"0000";
    tmp(81011) := x"0000";
    tmp(81012) := x"0000";
    tmp(81013) := x"0000";
    tmp(81014) := x"0000";
    tmp(81015) := x"0000";
    tmp(81016) := x"0000";
    tmp(81017) := x"0000";
    tmp(81018) := x"0000";
    tmp(81019) := x"0000";
    tmp(81020) := x"0000";
    tmp(81021) := x"0000";
    tmp(81022) := x"0000";
    tmp(81023) := x"0000";
    tmp(81024) := x"0000";
    tmp(81025) := x"0000";
    tmp(81026) := x"0000";
    tmp(81027) := x"0000";
    tmp(81028) := x"0000";
    tmp(81029) := x"0000";
    tmp(81030) := x"0000";
    tmp(81031) := x"0000";
    tmp(81032) := x"0000";
    tmp(81033) := x"0000";
    tmp(81034) := x"0000";
    tmp(81035) := x"0000";
    tmp(81036) := x"0000";
    tmp(81037) := x"0000";
    tmp(81038) := x"0000";
    tmp(81039) := x"0000";
    tmp(81040) := x"0000";
    tmp(81041) := x"0000";
    tmp(81042) := x"0000";
    tmp(81043) := x"0000";
    tmp(81044) := x"0000";
    tmp(81045) := x"0000";
    tmp(81046) := x"0000";
    tmp(81047) := x"0000";
    tmp(81048) := x"0000";
    tmp(81049) := x"0000";
    tmp(81050) := x"0000";
    tmp(81051) := x"0000";
    tmp(81052) := x"0000";
    tmp(81053) := x"0000";
    tmp(81054) := x"0000";
    tmp(81055) := x"0000";
    tmp(81056) := x"0000";
    tmp(81057) := x"0000";
    tmp(81058) := x"0000";
    tmp(81059) := x"0000";
    tmp(81060) := x"0000";
    tmp(81061) := x"0000";
    tmp(81062) := x"0000";
    tmp(81063) := x"0000";
    tmp(81064) := x"0000";
    tmp(81065) := x"0000";
    tmp(81066) := x"0000";
    tmp(81067) := x"0000";
    tmp(81068) := x"0000";
    tmp(81069) := x"0000";
    tmp(81070) := x"0000";
    tmp(81071) := x"0000";
    tmp(81072) := x"0000";
    tmp(81073) := x"0000";
    tmp(81074) := x"0000";
    tmp(81075) := x"0000";
    tmp(81076) := x"0000";
    tmp(81077) := x"0000";
    tmp(81078) := x"0000";
    tmp(81079) := x"0000";
    tmp(81080) := x"0000";
    tmp(81081) := x"0000";
    tmp(81082) := x"0000";
    tmp(81083) := x"0000";
    tmp(81084) := x"0000";
    tmp(81085) := x"0000";
    tmp(81086) := x"0000";
    tmp(81087) := x"0000";
    tmp(81088) := x"0000";
    tmp(81089) := x"0000";
    tmp(81090) := x"0000";
    tmp(81091) := x"0000";
    tmp(81092) := x"0000";
    tmp(81093) := x"0000";
    tmp(81094) := x"0000";
    tmp(81095) := x"0000";
    tmp(81096) := x"0000";
    tmp(81097) := x"0000";
    tmp(81098) := x"0000";
    tmp(81099) := x"0000";
    tmp(81100) := x"0000";
    tmp(81101) := x"0000";
    tmp(81102) := x"0000";
    tmp(81103) := x"0000";
    tmp(81104) := x"0000";
    tmp(81105) := x"0000";
    tmp(81106) := x"0000";
    tmp(81107) := x"0000";
    tmp(81108) := x"0000";
    tmp(81109) := x"0000";
    tmp(81110) := x"0000";
    tmp(81111) := x"0000";
    tmp(81112) := x"0000";
    tmp(81113) := x"0000";
    tmp(81114) := x"0000";
    tmp(81115) := x"0000";
    tmp(81116) := x"0000";
    tmp(81117) := x"0000";
    tmp(81118) := x"0000";
    tmp(81119) := x"0000";
    tmp(81120) := x"0000";
    tmp(81121) := x"0020";
    tmp(81122) := x"0020";
    tmp(81123) := x"0000";
    tmp(81124) := x"0000";
    tmp(81125) := x"0000";
    tmp(81126) := x"0000";
    tmp(81127) := x"0000";
    tmp(81128) := x"0000";
    tmp(81129) := x"0000";
    tmp(81130) := x"0000";
    tmp(81131) := x"0000";
    tmp(81132) := x"0000";
    tmp(81133) := x"0000";
    tmp(81134) := x"0000";
    tmp(81135) := x"0000";
    tmp(81136) := x"0000";
    tmp(81137) := x"0020";
    tmp(81138) := x"0020";
    tmp(81139) := x"0020";
    tmp(81140) := x"0020";
    tmp(81141) := x"0020";
    tmp(81142) := x"0020";
    tmp(81143) := x"0020";
    tmp(81144) := x"0020";
    tmp(81145) := x"0020";
    tmp(81146) := x"0020";
    tmp(81147) := x"0020";
    tmp(81148) := x"0020";
    tmp(81149) := x"0020";
    tmp(81150) := x"0020";
    tmp(81151) := x"0800";
    tmp(81152) := x"0000";
    tmp(81153) := x"0000";
    tmp(81154) := x"0800";
    tmp(81155) := x"0800";
    tmp(81156) := x"0800";
    tmp(81157) := x"0800";
    tmp(81158) := x"0800";
    tmp(81159) := x"0800";
    tmp(81160) := x"0800";
    tmp(81161) := x"0800";
    tmp(81162) := x"0800";
    tmp(81163) := x"0800";
    tmp(81164) := x"0800";
    tmp(81165) := x"0800";
    tmp(81166) := x"0800";
    tmp(81167) := x"0800";
    tmp(81168) := x"0800";
    tmp(81169) := x"0800";
    tmp(81170) := x"0800";
    tmp(81171) := x"0800";
    tmp(81172) := x"0800";
    tmp(81173) := x"0800";
    tmp(81174) := x"0800";
    tmp(81175) := x"1000";
    tmp(81176) := x"1000";
    tmp(81177) := x"1000";
    tmp(81178) := x"1000";
    tmp(81179) := x"0800";
    tmp(81180) := x"0800";
    tmp(81181) := x"0800";
    tmp(81182) := x"0800";
    tmp(81183) := x"0800";
    tmp(81184) := x"0800";
    tmp(81185) := x"0000";
    tmp(81186) := x"0000";
    tmp(81187) := x"0000";
    tmp(81188) := x"0000";
    tmp(81189) := x"0800";
    tmp(81190) := x"0800";
    tmp(81191) := x"0000";
    tmp(81192) := x"0000";
    tmp(81193) := x"0000";
    tmp(81194) := x"0800";
    tmp(81195) := x"1020";
    tmp(81196) := x"0000";
    tmp(81197) := x"0000";
    tmp(81198) := x"0000";
    tmp(81199) := x"0000";
    tmp(81200) := x"0800";
    tmp(81201) := x"0000";
    tmp(81202) := x"0000";
    tmp(81203) := x"0000";
    tmp(81204) := x"0000";
    tmp(81205) := x"0000";
    tmp(81206) := x"0800";
    tmp(81207) := x"1020";
    tmp(81208) := x"1020";
    tmp(81209) := x"0820";
    tmp(81210) := x"0800";
    tmp(81211) := x"0000";
    tmp(81212) := x"0000";
    tmp(81213) := x"0000";
    tmp(81214) := x"0000";
    tmp(81215) := x"0000";
    tmp(81216) := x"0000";
    tmp(81217) := x"0000";
    tmp(81218) := x"0000";
    tmp(81219) := x"0000";
    tmp(81220) := x"0000";
    tmp(81221) := x"0000";
    tmp(81222) := x"0000";
    tmp(81223) := x"0000";
    tmp(81224) := x"0000";
    tmp(81225) := x"0000";
    tmp(81226) := x"0000";
    tmp(81227) := x"0000";
    tmp(81228) := x"0000";
    tmp(81229) := x"0000";
    tmp(81230) := x"0000";
    tmp(81231) := x"0000";
    tmp(81232) := x"0000";
    tmp(81233) := x"0000";
    tmp(81234) := x"0000";
    tmp(81235) := x"0000";
    tmp(81236) := x"0000";
    tmp(81237) := x"0000";
    tmp(81238) := x"0000";
    tmp(81239) := x"0000";
    tmp(81240) := x"0000";
    tmp(81241) := x"0000";
    tmp(81242) := x"0000";
    tmp(81243) := x"0000";
    tmp(81244) := x"0000";
    tmp(81245) := x"0000";
    tmp(81246) := x"0000";
    tmp(81247) := x"0000";
    tmp(81248) := x"0000";
    tmp(81249) := x"0000";
    tmp(81250) := x"0000";
    tmp(81251) := x"0000";
    tmp(81252) := x"0000";
    tmp(81253) := x"0000";
    tmp(81254) := x"0000";
    tmp(81255) := x"0000";
    tmp(81256) := x"0000";
    tmp(81257) := x"0000";
    tmp(81258) := x"0000";
    tmp(81259) := x"0000";
    tmp(81260) := x"0000";
    tmp(81261) := x"0000";
    tmp(81262) := x"0000";
    tmp(81263) := x"0000";
    tmp(81264) := x"0000";
    tmp(81265) := x"0000";
    tmp(81266) := x"0000";
    tmp(81267) := x"0000";
    tmp(81268) := x"0000";
    tmp(81269) := x"0000";
    tmp(81270) := x"0000";
    tmp(81271) := x"0000";
    tmp(81272) := x"0000";
    tmp(81273) := x"0000";
    tmp(81274) := x"0000";
    tmp(81275) := x"0000";
    tmp(81276) := x"0000";
    tmp(81277) := x"0000";
    tmp(81278) := x"0000";
    tmp(81279) := x"0000";
    tmp(81280) := x"0000";
    tmp(81281) := x"0000";
    tmp(81282) := x"0000";
    tmp(81283) := x"0000";
    tmp(81284) := x"0000";
    tmp(81285) := x"0000";
    tmp(81286) := x"0000";
    tmp(81287) := x"0000";
    tmp(81288) := x"0000";
    tmp(81289) := x"0000";
    tmp(81290) := x"0000";
    tmp(81291) := x"0000";
    tmp(81292) := x"0000";
    tmp(81293) := x"0000";
    tmp(81294) := x"0000";
    tmp(81295) := x"0000";
    tmp(81296) := x"0000";
    tmp(81297) := x"0000";
    tmp(81298) := x"0000";
    tmp(81299) := x"0000";
    tmp(81300) := x"0000";
    tmp(81301) := x"0000";
    tmp(81302) := x"0000";
    tmp(81303) := x"0000";
    tmp(81304) := x"0000";
    tmp(81305) := x"0000";
    tmp(81306) := x"0000";
    tmp(81307) := x"0000";
    tmp(81308) := x"0000";
    tmp(81309) := x"0000";
    tmp(81310) := x"0000";
    tmp(81311) := x"0000";
    tmp(81312) := x"0000";
    tmp(81313) := x"0000";
    tmp(81314) := x"0000";
    tmp(81315) := x"0000";
    tmp(81316) := x"0000";
    tmp(81317) := x"0000";
    tmp(81318) := x"0000";
    tmp(81319) := x"0000";
    tmp(81320) := x"0000";
    tmp(81321) := x"0000";
    tmp(81322) := x"0000";
    tmp(81323) := x"0000";
    tmp(81324) := x"0000";
    tmp(81325) := x"0000";
    tmp(81326) := x"0000";
    tmp(81327) := x"0000";
    tmp(81328) := x"0000";
    tmp(81329) := x"0000";
    tmp(81330) := x"0000";
    tmp(81331) := x"0000";
    tmp(81332) := x"0000";
    tmp(81333) := x"0000";
    tmp(81334) := x"0000";
    tmp(81335) := x"0000";
    tmp(81336) := x"0000";
    tmp(81337) := x"0000";
    tmp(81338) := x"0000";
    tmp(81339) := x"0000";
    tmp(81340) := x"0000";
    tmp(81341) := x"0000";
    tmp(81342) := x"0000";
    tmp(81343) := x"0000";
    tmp(81344) := x"0000";
    tmp(81345) := x"0000";
    tmp(81346) := x"0000";
    tmp(81347) := x"0000";
    tmp(81348) := x"0000";
    tmp(81349) := x"0000";
    tmp(81350) := x"0000";
    tmp(81351) := x"0000";
    tmp(81352) := x"0000";
    tmp(81353) := x"0000";
    tmp(81354) := x"0000";
    tmp(81355) := x"0000";
    tmp(81356) := x"0000";
    tmp(81357) := x"0000";
    tmp(81358) := x"0000";
    tmp(81359) := x"0000";
    tmp(81360) := x"0000";
    tmp(81361) := x"0000";
    tmp(81362) := x"0020";
    tmp(81363) := x"0020";
    tmp(81364) := x"0020";
    tmp(81365) := x"0020";
    tmp(81366) := x"0020";
    tmp(81367) := x"0000";
    tmp(81368) := x"0000";
    tmp(81369) := x"0000";
    tmp(81370) := x"0000";
    tmp(81371) := x"0000";
    tmp(81372) := x"0000";
    tmp(81373) := x"0000";
    tmp(81374) := x"0000";
    tmp(81375) := x"0000";
    tmp(81376) := x"0020";
    tmp(81377) := x"0020";
    tmp(81378) := x"0020";
    tmp(81379) := x"0020";
    tmp(81380) := x"0020";
    tmp(81381) := x"0020";
    tmp(81382) := x"0020";
    tmp(81383) := x"0020";
    tmp(81384) := x"0020";
    tmp(81385) := x"0020";
    tmp(81386) := x"0020";
    tmp(81387) := x"0020";
    tmp(81388) := x"0020";
    tmp(81389) := x"0020";
    tmp(81390) := x"0820";
    tmp(81391) := x"0820";
    tmp(81392) := x"0800";
    tmp(81393) := x"0800";
    tmp(81394) := x"0800";
    tmp(81395) := x"0800";
    tmp(81396) := x"0800";
    tmp(81397) := x"0800";
    tmp(81398) := x"0800";
    tmp(81399) := x"0800";
    tmp(81400) := x"0800";
    tmp(81401) := x"0800";
    tmp(81402) := x"0800";
    tmp(81403) := x"0800";
    tmp(81404) := x"0800";
    tmp(81405) := x"0800";
    tmp(81406) := x"0800";
    tmp(81407) := x"0800";
    tmp(81408) := x"0800";
    tmp(81409) := x"0800";
    tmp(81410) := x"0800";
    tmp(81411) := x"0800";
    tmp(81412) := x"0800";
    tmp(81413) := x"0800";
    tmp(81414) := x"0800";
    tmp(81415) := x"0800";
    tmp(81416) := x"0800";
    tmp(81417) := x"0800";
    tmp(81418) := x"0800";
    tmp(81419) := x"0800";
    tmp(81420) := x"0800";
    tmp(81421) := x"0800";
    tmp(81422) := x"0800";
    tmp(81423) := x"0000";
    tmp(81424) := x"0000";
    tmp(81425) := x"0000";
    tmp(81426) := x"0800";
    tmp(81427) := x"0800";
    tmp(81428) := x"0800";
    tmp(81429) := x"0000";
    tmp(81430) := x"0000";
    tmp(81431) := x"0000";
    tmp(81432) := x"0000";
    tmp(81433) := x"1020";
    tmp(81434) := x"1000";
    tmp(81435) := x"0000";
    tmp(81436) := x"0000";
    tmp(81437) := x"0000";
    tmp(81438) := x"0000";
    tmp(81439) := x"0000";
    tmp(81440) := x"0000";
    tmp(81441) := x"0000";
    tmp(81442) := x"0000";
    tmp(81443) := x"0000";
    tmp(81444) := x"0800";
    tmp(81445) := x"1000";
    tmp(81446) := x"1020";
    tmp(81447) := x"1020";
    tmp(81448) := x"0800";
    tmp(81449) := x"0000";
    tmp(81450) := x"0000";
    tmp(81451) := x"0000";
    tmp(81452) := x"0000";
    tmp(81453) := x"0000";
    tmp(81454) := x"0000";
    tmp(81455) := x"0000";
    tmp(81456) := x"0000";
    tmp(81457) := x"0000";
    tmp(81458) := x"0000";
    tmp(81459) := x"0000";
    tmp(81460) := x"0000";
    tmp(81461) := x"0000";
    tmp(81462) := x"0000";
    tmp(81463) := x"0000";
    tmp(81464) := x"0000";
    tmp(81465) := x"0000";
    tmp(81466) := x"0000";
    tmp(81467) := x"0000";
    tmp(81468) := x"0000";
    tmp(81469) := x"0000";
    tmp(81470) := x"0000";
    tmp(81471) := x"0000";
    tmp(81472) := x"0000";
    tmp(81473) := x"0000";
    tmp(81474) := x"0000";
    tmp(81475) := x"0000";
    tmp(81476) := x"0000";
    tmp(81477) := x"0000";
    tmp(81478) := x"0000";
    tmp(81479) := x"0000";
    tmp(81480) := x"0000";
    tmp(81481) := x"0000";
    tmp(81482) := x"0000";
    tmp(81483) := x"0000";
    tmp(81484) := x"0000";
    tmp(81485) := x"0000";
    tmp(81486) := x"0000";
    tmp(81487) := x"0000";
    tmp(81488) := x"0000";
    tmp(81489) := x"0000";
    tmp(81490) := x"0000";
    tmp(81491) := x"0000";
    tmp(81492) := x"0000";
    tmp(81493) := x"0000";
    tmp(81494) := x"0000";
    tmp(81495) := x"0000";
    tmp(81496) := x"0000";
    tmp(81497) := x"0000";
    tmp(81498) := x"0000";
    tmp(81499) := x"0000";
    tmp(81500) := x"0000";
    tmp(81501) := x"0000";
    tmp(81502) := x"0000";
    tmp(81503) := x"0000";
    tmp(81504) := x"0000";
    tmp(81505) := x"0000";
    tmp(81506) := x"0000";
    tmp(81507) := x"0000";
    tmp(81508) := x"0000";
    tmp(81509) := x"0000";
    tmp(81510) := x"0000";
    tmp(81511) := x"0000";
    tmp(81512) := x"0000";
    tmp(81513) := x"0000";
    tmp(81514) := x"0000";
    tmp(81515) := x"0000";
    tmp(81516) := x"0000";
    tmp(81517) := x"0000";
    tmp(81518) := x"0000";
    tmp(81519) := x"0000";
    tmp(81520) := x"0000";
    tmp(81521) := x"0000";
    tmp(81522) := x"0000";
    tmp(81523) := x"0000";
    tmp(81524) := x"0000";
    tmp(81525) := x"0000";
    tmp(81526) := x"0000";
    tmp(81527) := x"0000";
    tmp(81528) := x"0000";
    tmp(81529) := x"0000";
    tmp(81530) := x"0000";
    tmp(81531) := x"0000";
    tmp(81532) := x"0000";
    tmp(81533) := x"0000";
    tmp(81534) := x"0000";
    tmp(81535) := x"0000";
    tmp(81536) := x"0000";
    tmp(81537) := x"0000";
    tmp(81538) := x"0000";
    tmp(81539) := x"0000";
    tmp(81540) := x"0000";
    tmp(81541) := x"0000";
    tmp(81542) := x"0000";
    tmp(81543) := x"0000";
    tmp(81544) := x"0000";
    tmp(81545) := x"0000";
    tmp(81546) := x"0000";
    tmp(81547) := x"0000";
    tmp(81548) := x"0000";
    tmp(81549) := x"0000";
    tmp(81550) := x"0000";
    tmp(81551) := x"0000";
    tmp(81552) := x"0000";
    tmp(81553) := x"0000";
    tmp(81554) := x"0000";
    tmp(81555) := x"0000";
    tmp(81556) := x"0000";
    tmp(81557) := x"0000";
    tmp(81558) := x"0000";
    tmp(81559) := x"0000";
    tmp(81560) := x"0000";
    tmp(81561) := x"0000";
    tmp(81562) := x"0000";
    tmp(81563) := x"0000";
    tmp(81564) := x"0000";
    tmp(81565) := x"0000";
    tmp(81566) := x"0000";
    tmp(81567) := x"0000";
    tmp(81568) := x"0000";
    tmp(81569) := x"0000";
    tmp(81570) := x"0000";
    tmp(81571) := x"0000";
    tmp(81572) := x"0000";
    tmp(81573) := x"0000";
    tmp(81574) := x"0000";
    tmp(81575) := x"0000";
    tmp(81576) := x"0000";
    tmp(81577) := x"0000";
    tmp(81578) := x"0000";
    tmp(81579) := x"0000";
    tmp(81580) := x"0000";
    tmp(81581) := x"0000";
    tmp(81582) := x"0000";
    tmp(81583) := x"0000";
    tmp(81584) := x"0000";
    tmp(81585) := x"0000";
    tmp(81586) := x"0000";
    tmp(81587) := x"0000";
    tmp(81588) := x"0000";
    tmp(81589) := x"0000";
    tmp(81590) := x"0000";
    tmp(81591) := x"0000";
    tmp(81592) := x"0000";
    tmp(81593) := x"0000";
    tmp(81594) := x"0000";
    tmp(81595) := x"0000";
    tmp(81596) := x"0000";
    tmp(81597) := x"0000";
    tmp(81598) := x"0000";
    tmp(81599) := x"0000";
    --end loop;
    return tmp;
  end init_rom;

  signal rom : memory_t := init_rom;

begin

  process(clk)
  begin
    if(rising_edge(clk)) then
      q <= rom(to_integer(unsigned(addr)));
    end if;
  end process;

end rtl;
---------------------------------------------------------------------------
